module Convo_Layer5#(
    parameter DATA_WIDHT = 32,
	parameter IMG_WIDHT = 44,
	parameter IMG_HEIGHT =44
)
(
    input [DATA_WIDHT*32-1:0] Data_In,
    input Valid_In,
    input clk,
    input rst,
    output [DATA_WIDHT*64-1:0] Data_Out,
    output Valid_Out
);
	wire[DATA_WIDHT*32-1:0] Data_Out_Kernel1, Data_Out_Kernel2, Data_Out_Kernel3, Data_Out_Kernel4, Data_Out_Kernel5, Data_Out_Kernel6, Data_Out_Kernel7, Data_Out_Kernel8, Data_Out_Kernel9, Data_Out_Kernel10, Data_Out_Kernel11, Data_Out_Kernel12, Data_Out_Kernel13, Data_Out_Kernel14, Data_Out_Kernel15, Data_Out_Kernel16, Data_Out_Kernel17, Data_Out_Kernel18, Data_Out_Kernel19, Data_Out_Kernel20, Data_Out_Kernel21, Data_Out_Kernel22, Data_Out_Kernel23, Data_Out_Kernel24, Data_Out_Kernel25, Data_Out_Kernel26, Data_Out_Kernel27, Data_Out_Kernel28, Data_Out_Kernel29, Data_Out_Kernel30, Data_Out_Kernel31, Data_Out_Kernel32, Data_Out_Kernel33, Data_Out_Kernel34, Data_Out_Kernel35, Data_Out_Kernel36, Data_Out_Kernel37, Data_Out_Kernel38, Data_Out_Kernel39, Data_Out_Kernel40, Data_Out_Kernel41, Data_Out_Kernel42, Data_Out_Kernel43, Data_Out_Kernel44, Data_Out_Kernel45, Data_Out_Kernel46, Data_Out_Kernel47, Data_Out_Kernel48, Data_Out_Kernel49, Data_Out_Kernel50, Data_Out_Kernel51, Data_Out_Kernel52, Data_Out_Kernel53, Data_Out_Kernel54, Data_Out_Kernel55, Data_Out_Kernel56, Data_Out_Kernel57, Data_Out_Kernel58, Data_Out_Kernel59, Data_Out_Kernel60, Data_Out_Kernel61, Data_Out_Kernel62, Data_Out_Kernel63, Data_Out_Kernel64;
	wire[31:0] add_k1_Data_Out, add_k2_Data_Out, add_k3_Data_Out, add_k4_Data_Out, add_k5_Data_Out, add_k6_Data_Out, add_k7_Data_Out, add_k8_Data_Out, add_k9_Data_Out, add_k10_Data_Out, add_k11_Data_Out, add_k12_Data_Out, add_k13_Data_Out, add_k14_Data_Out, add_k15_Data_Out, add_k16_Data_Out, add_k17_Data_Out, add_k18_Data_Out, add_k19_Data_Out, add_k20_Data_Out, add_k21_Data_Out, add_k22_Data_Out, add_k23_Data_Out, add_k24_Data_Out, add_k25_Data_Out, add_k26_Data_Out, add_k27_Data_Out, add_k28_Data_Out, add_k29_Data_Out, add_k30_Data_Out, add_k31_Data_Out, add_k32_Data_Out, add_k33_Data_Out, add_k34_Data_Out, add_k35_Data_Out, add_k36_Data_Out, add_k37_Data_Out, add_k38_Data_Out, add_k39_Data_Out, add_k40_Data_Out, add_k41_Data_Out, add_k42_Data_Out, add_k43_Data_Out, add_k44_Data_Out, add_k45_Data_Out, add_k46_Data_Out, add_k47_Data_Out, add_k48_Data_Out, add_k49_Data_Out, add_k50_Data_Out, add_k51_Data_Out, add_k52_Data_Out, add_k53_Data_Out, add_k54_Data_Out, add_k55_Data_Out, add_k56_Data_Out, add_k57_Data_Out, add_k58_Data_Out, add_k59_Data_Out, add_k60_Data_Out, add_k61_Data_Out, add_k62_Data_Out, add_k63_Data_Out, add_k64_Data_Out;

	wire add_kernel1_Valid_Out, add_kernel2_Valid_Out, add_kernel3_Valid_Out, add_kernel4_Valid_Out, add_kernel5_Valid_Out, add_kernel6_Valid_Out, add_kernel7_Valid_Out, add_kernel8_Valid_Out, add_kernel9_Valid_Out, add_kernel10_Valid_Out, add_kernel11_Valid_Out, add_kernel12_Valid_Out, add_kernel13_Valid_Out, add_kernel14_Valid_Out, add_kernel15_Valid_Out, add_kernel16_Valid_Out, add_kernel17_Valid_Out, add_kernel18_Valid_Out, add_kernel19_Valid_Out, add_kernel20_Valid_Out, add_kernel21_Valid_Out, add_kernel22_Valid_Out, add_kernel23_Valid_Out, add_kernel24_Valid_Out, add_kernel25_Valid_Out, add_kernel26_Valid_Out, add_kernel27_Valid_Out, add_kernel28_Valid_Out, add_kernel29_Valid_Out, add_kernel30_Valid_Out, add_kernel31_Valid_Out, add_kernel32_Valid_Out, add_kernel33_Valid_Out, add_kernel34_Valid_Out, add_kernel35_Valid_Out, add_kernel36_Valid_Out, add_kernel37_Valid_Out, add_kernel38_Valid_Out, add_kernel39_Valid_Out, add_kernel40_Valid_Out, add_kernel41_Valid_Out, add_kernel42_Valid_Out, add_kernel43_Valid_Out, add_kernel44_Valid_Out, add_kernel45_Valid_Out, add_kernel46_Valid_Out, add_kernel47_Valid_Out, add_kernel48_Valid_Out, add_kernel49_Valid_Out, add_kernel50_Valid_Out, add_kernel51_Valid_Out, add_kernel52_Valid_Out, add_kernel53_Valid_Out, add_kernel54_Valid_Out, add_kernel55_Valid_Out, add_kernel56_Valid_Out, add_kernel57_Valid_Out, add_kernel58_Valid_Out, add_kernel59_Valid_Out, add_kernel60_Valid_Out, add_kernel61_Valid_Out, add_kernel62_Valid_Out, add_kernel63_Valid_Out, add_kernel64_Valid_Out;

	wire channel1_Kernel1_Valid_Out, channel2_Kernel1_Valid_Out, channel3_Kernel1_Valid_Out, channel4_Kernel1_Valid_Out, channel5_Kernel1_Valid_Out, channel6_Kernel1_Valid_Out, channel7_Kernel1_Valid_Out, channel8_Kernel1_Valid_Out, channel9_Kernel1_Valid_Out, channel10_Kernel1_Valid_Out, channel11_Kernel1_Valid_Out, channel12_Kernel1_Valid_Out, channel13_Kernel1_Valid_Out, channel14_Kernel1_Valid_Out, channel15_Kernel1_Valid_Out, channel16_Kernel1_Valid_Out, channel17_Kernel1_Valid_Out, channel18_Kernel1_Valid_Out, channel19_Kernel1_Valid_Out, channel20_Kernel1_Valid_Out, channel21_Kernel1_Valid_Out, channel22_Kernel1_Valid_Out, channel23_Kernel1_Valid_Out, channel24_Kernel1_Valid_Out, channel25_Kernel1_Valid_Out, channel26_Kernel1_Valid_Out, channel27_Kernel1_Valid_Out, channel28_Kernel1_Valid_Out, channel29_Kernel1_Valid_Out, channel30_Kernel1_Valid_Out, channel31_Kernel1_Valid_Out, channel32_Kernel1_Valid_Out;

	assign add_kernel1=channel1_Kernel1_Valid_Out & channel2_Kernel1_Valid_Out & channel3_Kernel1_Valid_Out & channel4_Kernel1_Valid_Out & channel5_Kernel1_Valid_Out & channel6_Kernel1_Valid_Out & channel7_Kernel1_Valid_Out & channel8_Kernel1_Valid_Out & channel9_Kernel1_Valid_Out & channel10_Kernel1_Valid_Out & channel11_Kernel1_Valid_Out & channel12_Kernel1_Valid_Out & channel13_Kernel1_Valid_Out & channel14_Kernel1_Valid_Out & channel15_Kernel1_Valid_Out & channel16_Kernel1_Valid_Out & channel17_Kernel1_Valid_Out & channel18_Kernel1_Valid_Out & channel19_Kernel1_Valid_Out & channel20_Kernel1_Valid_Out & channel21_Kernel1_Valid_Out & channel22_Kernel1_Valid_Out & channel23_Kernel1_Valid_Out & channel24_Kernel1_Valid_Out & channel25_Kernel1_Valid_Out & channel26_Kernel1_Valid_Out & channel27_Kernel1_Valid_Out & channel28_Kernel1_Valid_Out & channel29_Kernel1_Valid_Out & channel30_Kernel1_Valid_Out & channel31_Kernel1_Valid_Out & channel32_Kernel1_Valid_Out;

	wire channel1_Kernel2_Valid_Out, channel2_Kernel2_Valid_Out, channel3_Kernel2_Valid_Out, channel4_Kernel2_Valid_Out, channel5_Kernel2_Valid_Out, channel6_Kernel2_Valid_Out, channel7_Kernel2_Valid_Out, channel8_Kernel2_Valid_Out, channel9_Kernel2_Valid_Out, channel10_Kernel2_Valid_Out, channel11_Kernel2_Valid_Out, channel12_Kernel2_Valid_Out, channel13_Kernel2_Valid_Out, channel14_Kernel2_Valid_Out, channel15_Kernel2_Valid_Out, channel16_Kernel2_Valid_Out, channel17_Kernel2_Valid_Out, channel18_Kernel2_Valid_Out, channel19_Kernel2_Valid_Out, channel20_Kernel2_Valid_Out, channel21_Kernel2_Valid_Out, channel22_Kernel2_Valid_Out, channel23_Kernel2_Valid_Out, channel24_Kernel2_Valid_Out, channel25_Kernel2_Valid_Out, channel26_Kernel2_Valid_Out, channel27_Kernel2_Valid_Out, channel28_Kernel2_Valid_Out, channel29_Kernel2_Valid_Out, channel30_Kernel2_Valid_Out, channel31_Kernel2_Valid_Out, channel32_Kernel2_Valid_Out;

	assign add_kernel2=channel1_Kernel2_Valid_Out & channel2_Kernel2_Valid_Out & channel3_Kernel2_Valid_Out & channel4_Kernel2_Valid_Out & channel5_Kernel2_Valid_Out & channel6_Kernel2_Valid_Out & channel7_Kernel2_Valid_Out & channel8_Kernel2_Valid_Out & channel9_Kernel2_Valid_Out & channel10_Kernel2_Valid_Out & channel11_Kernel2_Valid_Out & channel12_Kernel2_Valid_Out & channel13_Kernel2_Valid_Out & channel14_Kernel2_Valid_Out & channel15_Kernel2_Valid_Out & channel16_Kernel2_Valid_Out & channel17_Kernel2_Valid_Out & channel18_Kernel2_Valid_Out & channel19_Kernel2_Valid_Out & channel20_Kernel2_Valid_Out & channel21_Kernel2_Valid_Out & channel22_Kernel2_Valid_Out & channel23_Kernel2_Valid_Out & channel24_Kernel2_Valid_Out & channel25_Kernel2_Valid_Out & channel26_Kernel2_Valid_Out & channel27_Kernel2_Valid_Out & channel28_Kernel2_Valid_Out & channel29_Kernel2_Valid_Out & channel30_Kernel2_Valid_Out & channel31_Kernel2_Valid_Out & channel32_Kernel2_Valid_Out;

	wire channel1_Kernel3_Valid_Out, channel2_Kernel3_Valid_Out, channel3_Kernel3_Valid_Out, channel4_Kernel3_Valid_Out, channel5_Kernel3_Valid_Out, channel6_Kernel3_Valid_Out, channel7_Kernel3_Valid_Out, channel8_Kernel3_Valid_Out, channel9_Kernel3_Valid_Out, channel10_Kernel3_Valid_Out, channel11_Kernel3_Valid_Out, channel12_Kernel3_Valid_Out, channel13_Kernel3_Valid_Out, channel14_Kernel3_Valid_Out, channel15_Kernel3_Valid_Out, channel16_Kernel3_Valid_Out, channel17_Kernel3_Valid_Out, channel18_Kernel3_Valid_Out, channel19_Kernel3_Valid_Out, channel20_Kernel3_Valid_Out, channel21_Kernel3_Valid_Out, channel22_Kernel3_Valid_Out, channel23_Kernel3_Valid_Out, channel24_Kernel3_Valid_Out, channel25_Kernel3_Valid_Out, channel26_Kernel3_Valid_Out, channel27_Kernel3_Valid_Out, channel28_Kernel3_Valid_Out, channel29_Kernel3_Valid_Out, channel30_Kernel3_Valid_Out, channel31_Kernel3_Valid_Out, channel32_Kernel3_Valid_Out;

	assign add_kernel3=channel1_Kernel3_Valid_Out & channel2_Kernel3_Valid_Out & channel3_Kernel3_Valid_Out & channel4_Kernel3_Valid_Out & channel5_Kernel3_Valid_Out & channel6_Kernel3_Valid_Out & channel7_Kernel3_Valid_Out & channel8_Kernel3_Valid_Out & channel9_Kernel3_Valid_Out & channel10_Kernel3_Valid_Out & channel11_Kernel3_Valid_Out & channel12_Kernel3_Valid_Out & channel13_Kernel3_Valid_Out & channel14_Kernel3_Valid_Out & channel15_Kernel3_Valid_Out & channel16_Kernel3_Valid_Out & channel17_Kernel3_Valid_Out & channel18_Kernel3_Valid_Out & channel19_Kernel3_Valid_Out & channel20_Kernel3_Valid_Out & channel21_Kernel3_Valid_Out & channel22_Kernel3_Valid_Out & channel23_Kernel3_Valid_Out & channel24_Kernel3_Valid_Out & channel25_Kernel3_Valid_Out & channel26_Kernel3_Valid_Out & channel27_Kernel3_Valid_Out & channel28_Kernel3_Valid_Out & channel29_Kernel3_Valid_Out & channel30_Kernel3_Valid_Out & channel31_Kernel3_Valid_Out & channel32_Kernel3_Valid_Out;

	wire channel1_Kernel4_Valid_Out, channel2_Kernel4_Valid_Out, channel3_Kernel4_Valid_Out, channel4_Kernel4_Valid_Out, channel5_Kernel4_Valid_Out, channel6_Kernel4_Valid_Out, channel7_Kernel4_Valid_Out, channel8_Kernel4_Valid_Out, channel9_Kernel4_Valid_Out, channel10_Kernel4_Valid_Out, channel11_Kernel4_Valid_Out, channel12_Kernel4_Valid_Out, channel13_Kernel4_Valid_Out, channel14_Kernel4_Valid_Out, channel15_Kernel4_Valid_Out, channel16_Kernel4_Valid_Out, channel17_Kernel4_Valid_Out, channel18_Kernel4_Valid_Out, channel19_Kernel4_Valid_Out, channel20_Kernel4_Valid_Out, channel21_Kernel4_Valid_Out, channel22_Kernel4_Valid_Out, channel23_Kernel4_Valid_Out, channel24_Kernel4_Valid_Out, channel25_Kernel4_Valid_Out, channel26_Kernel4_Valid_Out, channel27_Kernel4_Valid_Out, channel28_Kernel4_Valid_Out, channel29_Kernel4_Valid_Out, channel30_Kernel4_Valid_Out, channel31_Kernel4_Valid_Out, channel32_Kernel4_Valid_Out;

	assign add_kernel4=channel1_Kernel4_Valid_Out & channel2_Kernel4_Valid_Out & channel3_Kernel4_Valid_Out & channel4_Kernel4_Valid_Out & channel5_Kernel4_Valid_Out & channel6_Kernel4_Valid_Out & channel7_Kernel4_Valid_Out & channel8_Kernel4_Valid_Out & channel9_Kernel4_Valid_Out & channel10_Kernel4_Valid_Out & channel11_Kernel4_Valid_Out & channel12_Kernel4_Valid_Out & channel13_Kernel4_Valid_Out & channel14_Kernel4_Valid_Out & channel15_Kernel4_Valid_Out & channel16_Kernel4_Valid_Out & channel17_Kernel4_Valid_Out & channel18_Kernel4_Valid_Out & channel19_Kernel4_Valid_Out & channel20_Kernel4_Valid_Out & channel21_Kernel4_Valid_Out & channel22_Kernel4_Valid_Out & channel23_Kernel4_Valid_Out & channel24_Kernel4_Valid_Out & channel25_Kernel4_Valid_Out & channel26_Kernel4_Valid_Out & channel27_Kernel4_Valid_Out & channel28_Kernel4_Valid_Out & channel29_Kernel4_Valid_Out & channel30_Kernel4_Valid_Out & channel31_Kernel4_Valid_Out & channel32_Kernel4_Valid_Out;

	wire channel1_Kernel5_Valid_Out, channel2_Kernel5_Valid_Out, channel3_Kernel5_Valid_Out, channel4_Kernel5_Valid_Out, channel5_Kernel5_Valid_Out, channel6_Kernel5_Valid_Out, channel7_Kernel5_Valid_Out, channel8_Kernel5_Valid_Out, channel9_Kernel5_Valid_Out, channel10_Kernel5_Valid_Out, channel11_Kernel5_Valid_Out, channel12_Kernel5_Valid_Out, channel13_Kernel5_Valid_Out, channel14_Kernel5_Valid_Out, channel15_Kernel5_Valid_Out, channel16_Kernel5_Valid_Out, channel17_Kernel5_Valid_Out, channel18_Kernel5_Valid_Out, channel19_Kernel5_Valid_Out, channel20_Kernel5_Valid_Out, channel21_Kernel5_Valid_Out, channel22_Kernel5_Valid_Out, channel23_Kernel5_Valid_Out, channel24_Kernel5_Valid_Out, channel25_Kernel5_Valid_Out, channel26_Kernel5_Valid_Out, channel27_Kernel5_Valid_Out, channel28_Kernel5_Valid_Out, channel29_Kernel5_Valid_Out, channel30_Kernel5_Valid_Out, channel31_Kernel5_Valid_Out, channel32_Kernel5_Valid_Out;

	assign add_kernel5=channel1_Kernel5_Valid_Out & channel2_Kernel5_Valid_Out & channel3_Kernel5_Valid_Out & channel4_Kernel5_Valid_Out & channel5_Kernel5_Valid_Out & channel6_Kernel5_Valid_Out & channel7_Kernel5_Valid_Out & channel8_Kernel5_Valid_Out & channel9_Kernel5_Valid_Out & channel10_Kernel5_Valid_Out & channel11_Kernel5_Valid_Out & channel12_Kernel5_Valid_Out & channel13_Kernel5_Valid_Out & channel14_Kernel5_Valid_Out & channel15_Kernel5_Valid_Out & channel16_Kernel5_Valid_Out & channel17_Kernel5_Valid_Out & channel18_Kernel5_Valid_Out & channel19_Kernel5_Valid_Out & channel20_Kernel5_Valid_Out & channel21_Kernel5_Valid_Out & channel22_Kernel5_Valid_Out & channel23_Kernel5_Valid_Out & channel24_Kernel5_Valid_Out & channel25_Kernel5_Valid_Out & channel26_Kernel5_Valid_Out & channel27_Kernel5_Valid_Out & channel28_Kernel5_Valid_Out & channel29_Kernel5_Valid_Out & channel30_Kernel5_Valid_Out & channel31_Kernel5_Valid_Out & channel32_Kernel5_Valid_Out;

	wire channel1_Kernel6_Valid_Out, channel2_Kernel6_Valid_Out, channel3_Kernel6_Valid_Out, channel4_Kernel6_Valid_Out, channel5_Kernel6_Valid_Out, channel6_Kernel6_Valid_Out, channel7_Kernel6_Valid_Out, channel8_Kernel6_Valid_Out, channel9_Kernel6_Valid_Out, channel10_Kernel6_Valid_Out, channel11_Kernel6_Valid_Out, channel12_Kernel6_Valid_Out, channel13_Kernel6_Valid_Out, channel14_Kernel6_Valid_Out, channel15_Kernel6_Valid_Out, channel16_Kernel6_Valid_Out, channel17_Kernel6_Valid_Out, channel18_Kernel6_Valid_Out, channel19_Kernel6_Valid_Out, channel20_Kernel6_Valid_Out, channel21_Kernel6_Valid_Out, channel22_Kernel6_Valid_Out, channel23_Kernel6_Valid_Out, channel24_Kernel6_Valid_Out, channel25_Kernel6_Valid_Out, channel26_Kernel6_Valid_Out, channel27_Kernel6_Valid_Out, channel28_Kernel6_Valid_Out, channel29_Kernel6_Valid_Out, channel30_Kernel6_Valid_Out, channel31_Kernel6_Valid_Out, channel32_Kernel6_Valid_Out;

	assign add_kernel6=channel1_Kernel6_Valid_Out & channel2_Kernel6_Valid_Out & channel3_Kernel6_Valid_Out & channel4_Kernel6_Valid_Out & channel5_Kernel6_Valid_Out & channel6_Kernel6_Valid_Out & channel7_Kernel6_Valid_Out & channel8_Kernel6_Valid_Out & channel9_Kernel6_Valid_Out & channel10_Kernel6_Valid_Out & channel11_Kernel6_Valid_Out & channel12_Kernel6_Valid_Out & channel13_Kernel6_Valid_Out & channel14_Kernel6_Valid_Out & channel15_Kernel6_Valid_Out & channel16_Kernel6_Valid_Out & channel17_Kernel6_Valid_Out & channel18_Kernel6_Valid_Out & channel19_Kernel6_Valid_Out & channel20_Kernel6_Valid_Out & channel21_Kernel6_Valid_Out & channel22_Kernel6_Valid_Out & channel23_Kernel6_Valid_Out & channel24_Kernel6_Valid_Out & channel25_Kernel6_Valid_Out & channel26_Kernel6_Valid_Out & channel27_Kernel6_Valid_Out & channel28_Kernel6_Valid_Out & channel29_Kernel6_Valid_Out & channel30_Kernel6_Valid_Out & channel31_Kernel6_Valid_Out & channel32_Kernel6_Valid_Out;

	wire channel1_Kernel7_Valid_Out, channel2_Kernel7_Valid_Out, channel3_Kernel7_Valid_Out, channel4_Kernel7_Valid_Out, channel5_Kernel7_Valid_Out, channel6_Kernel7_Valid_Out, channel7_Kernel7_Valid_Out, channel8_Kernel7_Valid_Out, channel9_Kernel7_Valid_Out, channel10_Kernel7_Valid_Out, channel11_Kernel7_Valid_Out, channel12_Kernel7_Valid_Out, channel13_Kernel7_Valid_Out, channel14_Kernel7_Valid_Out, channel15_Kernel7_Valid_Out, channel16_Kernel7_Valid_Out, channel17_Kernel7_Valid_Out, channel18_Kernel7_Valid_Out, channel19_Kernel7_Valid_Out, channel20_Kernel7_Valid_Out, channel21_Kernel7_Valid_Out, channel22_Kernel7_Valid_Out, channel23_Kernel7_Valid_Out, channel24_Kernel7_Valid_Out, channel25_Kernel7_Valid_Out, channel26_Kernel7_Valid_Out, channel27_Kernel7_Valid_Out, channel28_Kernel7_Valid_Out, channel29_Kernel7_Valid_Out, channel30_Kernel7_Valid_Out, channel31_Kernel7_Valid_Out, channel32_Kernel7_Valid_Out;

	assign add_kernel7=channel1_Kernel7_Valid_Out & channel2_Kernel7_Valid_Out & channel3_Kernel7_Valid_Out & channel4_Kernel7_Valid_Out & channel5_Kernel7_Valid_Out & channel6_Kernel7_Valid_Out & channel7_Kernel7_Valid_Out & channel8_Kernel7_Valid_Out & channel9_Kernel7_Valid_Out & channel10_Kernel7_Valid_Out & channel11_Kernel7_Valid_Out & channel12_Kernel7_Valid_Out & channel13_Kernel7_Valid_Out & channel14_Kernel7_Valid_Out & channel15_Kernel7_Valid_Out & channel16_Kernel7_Valid_Out & channel17_Kernel7_Valid_Out & channel18_Kernel7_Valid_Out & channel19_Kernel7_Valid_Out & channel20_Kernel7_Valid_Out & channel21_Kernel7_Valid_Out & channel22_Kernel7_Valid_Out & channel23_Kernel7_Valid_Out & channel24_Kernel7_Valid_Out & channel25_Kernel7_Valid_Out & channel26_Kernel7_Valid_Out & channel27_Kernel7_Valid_Out & channel28_Kernel7_Valid_Out & channel29_Kernel7_Valid_Out & channel30_Kernel7_Valid_Out & channel31_Kernel7_Valid_Out & channel32_Kernel7_Valid_Out;

	wire channel1_Kernel8_Valid_Out, channel2_Kernel8_Valid_Out, channel3_Kernel8_Valid_Out, channel4_Kernel8_Valid_Out, channel5_Kernel8_Valid_Out, channel6_Kernel8_Valid_Out, channel7_Kernel8_Valid_Out, channel8_Kernel8_Valid_Out, channel9_Kernel8_Valid_Out, channel10_Kernel8_Valid_Out, channel11_Kernel8_Valid_Out, channel12_Kernel8_Valid_Out, channel13_Kernel8_Valid_Out, channel14_Kernel8_Valid_Out, channel15_Kernel8_Valid_Out, channel16_Kernel8_Valid_Out, channel17_Kernel8_Valid_Out, channel18_Kernel8_Valid_Out, channel19_Kernel8_Valid_Out, channel20_Kernel8_Valid_Out, channel21_Kernel8_Valid_Out, channel22_Kernel8_Valid_Out, channel23_Kernel8_Valid_Out, channel24_Kernel8_Valid_Out, channel25_Kernel8_Valid_Out, channel26_Kernel8_Valid_Out, channel27_Kernel8_Valid_Out, channel28_Kernel8_Valid_Out, channel29_Kernel8_Valid_Out, channel30_Kernel8_Valid_Out, channel31_Kernel8_Valid_Out, channel32_Kernel8_Valid_Out;

	assign add_kernel8=channel1_Kernel8_Valid_Out & channel2_Kernel8_Valid_Out & channel3_Kernel8_Valid_Out & channel4_Kernel8_Valid_Out & channel5_Kernel8_Valid_Out & channel6_Kernel8_Valid_Out & channel7_Kernel8_Valid_Out & channel8_Kernel8_Valid_Out & channel9_Kernel8_Valid_Out & channel10_Kernel8_Valid_Out & channel11_Kernel8_Valid_Out & channel12_Kernel8_Valid_Out & channel13_Kernel8_Valid_Out & channel14_Kernel8_Valid_Out & channel15_Kernel8_Valid_Out & channel16_Kernel8_Valid_Out & channel17_Kernel8_Valid_Out & channel18_Kernel8_Valid_Out & channel19_Kernel8_Valid_Out & channel20_Kernel8_Valid_Out & channel21_Kernel8_Valid_Out & channel22_Kernel8_Valid_Out & channel23_Kernel8_Valid_Out & channel24_Kernel8_Valid_Out & channel25_Kernel8_Valid_Out & channel26_Kernel8_Valid_Out & channel27_Kernel8_Valid_Out & channel28_Kernel8_Valid_Out & channel29_Kernel8_Valid_Out & channel30_Kernel8_Valid_Out & channel31_Kernel8_Valid_Out & channel32_Kernel8_Valid_Out;

	wire channel1_Kernel9_Valid_Out, channel2_Kernel9_Valid_Out, channel3_Kernel9_Valid_Out, channel4_Kernel9_Valid_Out, channel5_Kernel9_Valid_Out, channel6_Kernel9_Valid_Out, channel7_Kernel9_Valid_Out, channel8_Kernel9_Valid_Out, channel9_Kernel9_Valid_Out, channel10_Kernel9_Valid_Out, channel11_Kernel9_Valid_Out, channel12_Kernel9_Valid_Out, channel13_Kernel9_Valid_Out, channel14_Kernel9_Valid_Out, channel15_Kernel9_Valid_Out, channel16_Kernel9_Valid_Out, channel17_Kernel9_Valid_Out, channel18_Kernel9_Valid_Out, channel19_Kernel9_Valid_Out, channel20_Kernel9_Valid_Out, channel21_Kernel9_Valid_Out, channel22_Kernel9_Valid_Out, channel23_Kernel9_Valid_Out, channel24_Kernel9_Valid_Out, channel25_Kernel9_Valid_Out, channel26_Kernel9_Valid_Out, channel27_Kernel9_Valid_Out, channel28_Kernel9_Valid_Out, channel29_Kernel9_Valid_Out, channel30_Kernel9_Valid_Out, channel31_Kernel9_Valid_Out, channel32_Kernel9_Valid_Out;

	assign add_kernel9=channel1_Kernel9_Valid_Out & channel2_Kernel9_Valid_Out & channel3_Kernel9_Valid_Out & channel4_Kernel9_Valid_Out & channel5_Kernel9_Valid_Out & channel6_Kernel9_Valid_Out & channel7_Kernel9_Valid_Out & channel8_Kernel9_Valid_Out & channel9_Kernel9_Valid_Out & channel10_Kernel9_Valid_Out & channel11_Kernel9_Valid_Out & channel12_Kernel9_Valid_Out & channel13_Kernel9_Valid_Out & channel14_Kernel9_Valid_Out & channel15_Kernel9_Valid_Out & channel16_Kernel9_Valid_Out & channel17_Kernel9_Valid_Out & channel18_Kernel9_Valid_Out & channel19_Kernel9_Valid_Out & channel20_Kernel9_Valid_Out & channel21_Kernel9_Valid_Out & channel22_Kernel9_Valid_Out & channel23_Kernel9_Valid_Out & channel24_Kernel9_Valid_Out & channel25_Kernel9_Valid_Out & channel26_Kernel9_Valid_Out & channel27_Kernel9_Valid_Out & channel28_Kernel9_Valid_Out & channel29_Kernel9_Valid_Out & channel30_Kernel9_Valid_Out & channel31_Kernel9_Valid_Out & channel32_Kernel9_Valid_Out;

	wire channel1_Kernel10_Valid_Out, channel2_Kernel10_Valid_Out, channel3_Kernel10_Valid_Out, channel4_Kernel10_Valid_Out, channel5_Kernel10_Valid_Out, channel6_Kernel10_Valid_Out, channel7_Kernel10_Valid_Out, channel8_Kernel10_Valid_Out, channel9_Kernel10_Valid_Out, channel10_Kernel10_Valid_Out, channel11_Kernel10_Valid_Out, channel12_Kernel10_Valid_Out, channel13_Kernel10_Valid_Out, channel14_Kernel10_Valid_Out, channel15_Kernel10_Valid_Out, channel16_Kernel10_Valid_Out, channel17_Kernel10_Valid_Out, channel18_Kernel10_Valid_Out, channel19_Kernel10_Valid_Out, channel20_Kernel10_Valid_Out, channel21_Kernel10_Valid_Out, channel22_Kernel10_Valid_Out, channel23_Kernel10_Valid_Out, channel24_Kernel10_Valid_Out, channel25_Kernel10_Valid_Out, channel26_Kernel10_Valid_Out, channel27_Kernel10_Valid_Out, channel28_Kernel10_Valid_Out, channel29_Kernel10_Valid_Out, channel30_Kernel10_Valid_Out, channel31_Kernel10_Valid_Out, channel32_Kernel10_Valid_Out;

	assign add_kernel10=channel1_Kernel10_Valid_Out & channel2_Kernel10_Valid_Out & channel3_Kernel10_Valid_Out & channel4_Kernel10_Valid_Out & channel5_Kernel10_Valid_Out & channel6_Kernel10_Valid_Out & channel7_Kernel10_Valid_Out & channel8_Kernel10_Valid_Out & channel9_Kernel10_Valid_Out & channel10_Kernel10_Valid_Out & channel11_Kernel10_Valid_Out & channel12_Kernel10_Valid_Out & channel13_Kernel10_Valid_Out & channel14_Kernel10_Valid_Out & channel15_Kernel10_Valid_Out & channel16_Kernel10_Valid_Out & channel17_Kernel10_Valid_Out & channel18_Kernel10_Valid_Out & channel19_Kernel10_Valid_Out & channel20_Kernel10_Valid_Out & channel21_Kernel10_Valid_Out & channel22_Kernel10_Valid_Out & channel23_Kernel10_Valid_Out & channel24_Kernel10_Valid_Out & channel25_Kernel10_Valid_Out & channel26_Kernel10_Valid_Out & channel27_Kernel10_Valid_Out & channel28_Kernel10_Valid_Out & channel29_Kernel10_Valid_Out & channel30_Kernel10_Valid_Out & channel31_Kernel10_Valid_Out & channel32_Kernel10_Valid_Out;

	wire channel1_Kernel11_Valid_Out, channel2_Kernel11_Valid_Out, channel3_Kernel11_Valid_Out, channel4_Kernel11_Valid_Out, channel5_Kernel11_Valid_Out, channel6_Kernel11_Valid_Out, channel7_Kernel11_Valid_Out, channel8_Kernel11_Valid_Out, channel9_Kernel11_Valid_Out, channel10_Kernel11_Valid_Out, channel11_Kernel11_Valid_Out, channel12_Kernel11_Valid_Out, channel13_Kernel11_Valid_Out, channel14_Kernel11_Valid_Out, channel15_Kernel11_Valid_Out, channel16_Kernel11_Valid_Out, channel17_Kernel11_Valid_Out, channel18_Kernel11_Valid_Out, channel19_Kernel11_Valid_Out, channel20_Kernel11_Valid_Out, channel21_Kernel11_Valid_Out, channel22_Kernel11_Valid_Out, channel23_Kernel11_Valid_Out, channel24_Kernel11_Valid_Out, channel25_Kernel11_Valid_Out, channel26_Kernel11_Valid_Out, channel27_Kernel11_Valid_Out, channel28_Kernel11_Valid_Out, channel29_Kernel11_Valid_Out, channel30_Kernel11_Valid_Out, channel31_Kernel11_Valid_Out, channel32_Kernel11_Valid_Out;

	assign add_kernel11=channel1_Kernel11_Valid_Out & channel2_Kernel11_Valid_Out & channel3_Kernel11_Valid_Out & channel4_Kernel11_Valid_Out & channel5_Kernel11_Valid_Out & channel6_Kernel11_Valid_Out & channel7_Kernel11_Valid_Out & channel8_Kernel11_Valid_Out & channel9_Kernel11_Valid_Out & channel10_Kernel11_Valid_Out & channel11_Kernel11_Valid_Out & channel12_Kernel11_Valid_Out & channel13_Kernel11_Valid_Out & channel14_Kernel11_Valid_Out & channel15_Kernel11_Valid_Out & channel16_Kernel11_Valid_Out & channel17_Kernel11_Valid_Out & channel18_Kernel11_Valid_Out & channel19_Kernel11_Valid_Out & channel20_Kernel11_Valid_Out & channel21_Kernel11_Valid_Out & channel22_Kernel11_Valid_Out & channel23_Kernel11_Valid_Out & channel24_Kernel11_Valid_Out & channel25_Kernel11_Valid_Out & channel26_Kernel11_Valid_Out & channel27_Kernel11_Valid_Out & channel28_Kernel11_Valid_Out & channel29_Kernel11_Valid_Out & channel30_Kernel11_Valid_Out & channel31_Kernel11_Valid_Out & channel32_Kernel11_Valid_Out;

	wire channel1_Kernel12_Valid_Out, channel2_Kernel12_Valid_Out, channel3_Kernel12_Valid_Out, channel4_Kernel12_Valid_Out, channel5_Kernel12_Valid_Out, channel6_Kernel12_Valid_Out, channel7_Kernel12_Valid_Out, channel8_Kernel12_Valid_Out, channel9_Kernel12_Valid_Out, channel10_Kernel12_Valid_Out, channel11_Kernel12_Valid_Out, channel12_Kernel12_Valid_Out, channel13_Kernel12_Valid_Out, channel14_Kernel12_Valid_Out, channel15_Kernel12_Valid_Out, channel16_Kernel12_Valid_Out, channel17_Kernel12_Valid_Out, channel18_Kernel12_Valid_Out, channel19_Kernel12_Valid_Out, channel20_Kernel12_Valid_Out, channel21_Kernel12_Valid_Out, channel22_Kernel12_Valid_Out, channel23_Kernel12_Valid_Out, channel24_Kernel12_Valid_Out, channel25_Kernel12_Valid_Out, channel26_Kernel12_Valid_Out, channel27_Kernel12_Valid_Out, channel28_Kernel12_Valid_Out, channel29_Kernel12_Valid_Out, channel30_Kernel12_Valid_Out, channel31_Kernel12_Valid_Out, channel32_Kernel12_Valid_Out;

	assign add_kernel12=channel1_Kernel12_Valid_Out & channel2_Kernel12_Valid_Out & channel3_Kernel12_Valid_Out & channel4_Kernel12_Valid_Out & channel5_Kernel12_Valid_Out & channel6_Kernel12_Valid_Out & channel7_Kernel12_Valid_Out & channel8_Kernel12_Valid_Out & channel9_Kernel12_Valid_Out & channel10_Kernel12_Valid_Out & channel11_Kernel12_Valid_Out & channel12_Kernel12_Valid_Out & channel13_Kernel12_Valid_Out & channel14_Kernel12_Valid_Out & channel15_Kernel12_Valid_Out & channel16_Kernel12_Valid_Out & channel17_Kernel12_Valid_Out & channel18_Kernel12_Valid_Out & channel19_Kernel12_Valid_Out & channel20_Kernel12_Valid_Out & channel21_Kernel12_Valid_Out & channel22_Kernel12_Valid_Out & channel23_Kernel12_Valid_Out & channel24_Kernel12_Valid_Out & channel25_Kernel12_Valid_Out & channel26_Kernel12_Valid_Out & channel27_Kernel12_Valid_Out & channel28_Kernel12_Valid_Out & channel29_Kernel12_Valid_Out & channel30_Kernel12_Valid_Out & channel31_Kernel12_Valid_Out & channel32_Kernel12_Valid_Out;

	wire channel1_Kernel13_Valid_Out, channel2_Kernel13_Valid_Out, channel3_Kernel13_Valid_Out, channel4_Kernel13_Valid_Out, channel5_Kernel13_Valid_Out, channel6_Kernel13_Valid_Out, channel7_Kernel13_Valid_Out, channel8_Kernel13_Valid_Out, channel9_Kernel13_Valid_Out, channel10_Kernel13_Valid_Out, channel11_Kernel13_Valid_Out, channel12_Kernel13_Valid_Out, channel13_Kernel13_Valid_Out, channel14_Kernel13_Valid_Out, channel15_Kernel13_Valid_Out, channel16_Kernel13_Valid_Out, channel17_Kernel13_Valid_Out, channel18_Kernel13_Valid_Out, channel19_Kernel13_Valid_Out, channel20_Kernel13_Valid_Out, channel21_Kernel13_Valid_Out, channel22_Kernel13_Valid_Out, channel23_Kernel13_Valid_Out, channel24_Kernel13_Valid_Out, channel25_Kernel13_Valid_Out, channel26_Kernel13_Valid_Out, channel27_Kernel13_Valid_Out, channel28_Kernel13_Valid_Out, channel29_Kernel13_Valid_Out, channel30_Kernel13_Valid_Out, channel31_Kernel13_Valid_Out, channel32_Kernel13_Valid_Out;

	assign add_kernel13=channel1_Kernel13_Valid_Out & channel2_Kernel13_Valid_Out & channel3_Kernel13_Valid_Out & channel4_Kernel13_Valid_Out & channel5_Kernel13_Valid_Out & channel6_Kernel13_Valid_Out & channel7_Kernel13_Valid_Out & channel8_Kernel13_Valid_Out & channel9_Kernel13_Valid_Out & channel10_Kernel13_Valid_Out & channel11_Kernel13_Valid_Out & channel12_Kernel13_Valid_Out & channel13_Kernel13_Valid_Out & channel14_Kernel13_Valid_Out & channel15_Kernel13_Valid_Out & channel16_Kernel13_Valid_Out & channel17_Kernel13_Valid_Out & channel18_Kernel13_Valid_Out & channel19_Kernel13_Valid_Out & channel20_Kernel13_Valid_Out & channel21_Kernel13_Valid_Out & channel22_Kernel13_Valid_Out & channel23_Kernel13_Valid_Out & channel24_Kernel13_Valid_Out & channel25_Kernel13_Valid_Out & channel26_Kernel13_Valid_Out & channel27_Kernel13_Valid_Out & channel28_Kernel13_Valid_Out & channel29_Kernel13_Valid_Out & channel30_Kernel13_Valid_Out & channel31_Kernel13_Valid_Out & channel32_Kernel13_Valid_Out;

	wire channel1_Kernel14_Valid_Out, channel2_Kernel14_Valid_Out, channel3_Kernel14_Valid_Out, channel4_Kernel14_Valid_Out, channel5_Kernel14_Valid_Out, channel6_Kernel14_Valid_Out, channel7_Kernel14_Valid_Out, channel8_Kernel14_Valid_Out, channel9_Kernel14_Valid_Out, channel10_Kernel14_Valid_Out, channel11_Kernel14_Valid_Out, channel12_Kernel14_Valid_Out, channel13_Kernel14_Valid_Out, channel14_Kernel14_Valid_Out, channel15_Kernel14_Valid_Out, channel16_Kernel14_Valid_Out, channel17_Kernel14_Valid_Out, channel18_Kernel14_Valid_Out, channel19_Kernel14_Valid_Out, channel20_Kernel14_Valid_Out, channel21_Kernel14_Valid_Out, channel22_Kernel14_Valid_Out, channel23_Kernel14_Valid_Out, channel24_Kernel14_Valid_Out, channel25_Kernel14_Valid_Out, channel26_Kernel14_Valid_Out, channel27_Kernel14_Valid_Out, channel28_Kernel14_Valid_Out, channel29_Kernel14_Valid_Out, channel30_Kernel14_Valid_Out, channel31_Kernel14_Valid_Out, channel32_Kernel14_Valid_Out;

	assign add_kernel14=channel1_Kernel14_Valid_Out & channel2_Kernel14_Valid_Out & channel3_Kernel14_Valid_Out & channel4_Kernel14_Valid_Out & channel5_Kernel14_Valid_Out & channel6_Kernel14_Valid_Out & channel7_Kernel14_Valid_Out & channel8_Kernel14_Valid_Out & channel9_Kernel14_Valid_Out & channel10_Kernel14_Valid_Out & channel11_Kernel14_Valid_Out & channel12_Kernel14_Valid_Out & channel13_Kernel14_Valid_Out & channel14_Kernel14_Valid_Out & channel15_Kernel14_Valid_Out & channel16_Kernel14_Valid_Out & channel17_Kernel14_Valid_Out & channel18_Kernel14_Valid_Out & channel19_Kernel14_Valid_Out & channel20_Kernel14_Valid_Out & channel21_Kernel14_Valid_Out & channel22_Kernel14_Valid_Out & channel23_Kernel14_Valid_Out & channel24_Kernel14_Valid_Out & channel25_Kernel14_Valid_Out & channel26_Kernel14_Valid_Out & channel27_Kernel14_Valid_Out & channel28_Kernel14_Valid_Out & channel29_Kernel14_Valid_Out & channel30_Kernel14_Valid_Out & channel31_Kernel14_Valid_Out & channel32_Kernel14_Valid_Out;

	wire channel1_Kernel15_Valid_Out, channel2_Kernel15_Valid_Out, channel3_Kernel15_Valid_Out, channel4_Kernel15_Valid_Out, channel5_Kernel15_Valid_Out, channel6_Kernel15_Valid_Out, channel7_Kernel15_Valid_Out, channel8_Kernel15_Valid_Out, channel9_Kernel15_Valid_Out, channel10_Kernel15_Valid_Out, channel11_Kernel15_Valid_Out, channel12_Kernel15_Valid_Out, channel13_Kernel15_Valid_Out, channel14_Kernel15_Valid_Out, channel15_Kernel15_Valid_Out, channel16_Kernel15_Valid_Out, channel17_Kernel15_Valid_Out, channel18_Kernel15_Valid_Out, channel19_Kernel15_Valid_Out, channel20_Kernel15_Valid_Out, channel21_Kernel15_Valid_Out, channel22_Kernel15_Valid_Out, channel23_Kernel15_Valid_Out, channel24_Kernel15_Valid_Out, channel25_Kernel15_Valid_Out, channel26_Kernel15_Valid_Out, channel27_Kernel15_Valid_Out, channel28_Kernel15_Valid_Out, channel29_Kernel15_Valid_Out, channel30_Kernel15_Valid_Out, channel31_Kernel15_Valid_Out, channel32_Kernel15_Valid_Out;

	assign add_kernel15=channel1_Kernel15_Valid_Out & channel2_Kernel15_Valid_Out & channel3_Kernel15_Valid_Out & channel4_Kernel15_Valid_Out & channel5_Kernel15_Valid_Out & channel6_Kernel15_Valid_Out & channel7_Kernel15_Valid_Out & channel8_Kernel15_Valid_Out & channel9_Kernel15_Valid_Out & channel10_Kernel15_Valid_Out & channel11_Kernel15_Valid_Out & channel12_Kernel15_Valid_Out & channel13_Kernel15_Valid_Out & channel14_Kernel15_Valid_Out & channel15_Kernel15_Valid_Out & channel16_Kernel15_Valid_Out & channel17_Kernel15_Valid_Out & channel18_Kernel15_Valid_Out & channel19_Kernel15_Valid_Out & channel20_Kernel15_Valid_Out & channel21_Kernel15_Valid_Out & channel22_Kernel15_Valid_Out & channel23_Kernel15_Valid_Out & channel24_Kernel15_Valid_Out & channel25_Kernel15_Valid_Out & channel26_Kernel15_Valid_Out & channel27_Kernel15_Valid_Out & channel28_Kernel15_Valid_Out & channel29_Kernel15_Valid_Out & channel30_Kernel15_Valid_Out & channel31_Kernel15_Valid_Out & channel32_Kernel15_Valid_Out;

	wire channel1_Kernel16_Valid_Out, channel2_Kernel16_Valid_Out, channel3_Kernel16_Valid_Out, channel4_Kernel16_Valid_Out, channel5_Kernel16_Valid_Out, channel6_Kernel16_Valid_Out, channel7_Kernel16_Valid_Out, channel8_Kernel16_Valid_Out, channel9_Kernel16_Valid_Out, channel10_Kernel16_Valid_Out, channel11_Kernel16_Valid_Out, channel12_Kernel16_Valid_Out, channel13_Kernel16_Valid_Out, channel14_Kernel16_Valid_Out, channel15_Kernel16_Valid_Out, channel16_Kernel16_Valid_Out, channel17_Kernel16_Valid_Out, channel18_Kernel16_Valid_Out, channel19_Kernel16_Valid_Out, channel20_Kernel16_Valid_Out, channel21_Kernel16_Valid_Out, channel22_Kernel16_Valid_Out, channel23_Kernel16_Valid_Out, channel24_Kernel16_Valid_Out, channel25_Kernel16_Valid_Out, channel26_Kernel16_Valid_Out, channel27_Kernel16_Valid_Out, channel28_Kernel16_Valid_Out, channel29_Kernel16_Valid_Out, channel30_Kernel16_Valid_Out, channel31_Kernel16_Valid_Out, channel32_Kernel16_Valid_Out;

	assign add_kernel16=channel1_Kernel16_Valid_Out & channel2_Kernel16_Valid_Out & channel3_Kernel16_Valid_Out & channel4_Kernel16_Valid_Out & channel5_Kernel16_Valid_Out & channel6_Kernel16_Valid_Out & channel7_Kernel16_Valid_Out & channel8_Kernel16_Valid_Out & channel9_Kernel16_Valid_Out & channel10_Kernel16_Valid_Out & channel11_Kernel16_Valid_Out & channel12_Kernel16_Valid_Out & channel13_Kernel16_Valid_Out & channel14_Kernel16_Valid_Out & channel15_Kernel16_Valid_Out & channel16_Kernel16_Valid_Out & channel17_Kernel16_Valid_Out & channel18_Kernel16_Valid_Out & channel19_Kernel16_Valid_Out & channel20_Kernel16_Valid_Out & channel21_Kernel16_Valid_Out & channel22_Kernel16_Valid_Out & channel23_Kernel16_Valid_Out & channel24_Kernel16_Valid_Out & channel25_Kernel16_Valid_Out & channel26_Kernel16_Valid_Out & channel27_Kernel16_Valid_Out & channel28_Kernel16_Valid_Out & channel29_Kernel16_Valid_Out & channel30_Kernel16_Valid_Out & channel31_Kernel16_Valid_Out & channel32_Kernel16_Valid_Out;

	wire channel1_Kernel17_Valid_Out, channel2_Kernel17_Valid_Out, channel3_Kernel17_Valid_Out, channel4_Kernel17_Valid_Out, channel5_Kernel17_Valid_Out, channel6_Kernel17_Valid_Out, channel7_Kernel17_Valid_Out, channel8_Kernel17_Valid_Out, channel9_Kernel17_Valid_Out, channel10_Kernel17_Valid_Out, channel11_Kernel17_Valid_Out, channel12_Kernel17_Valid_Out, channel13_Kernel17_Valid_Out, channel14_Kernel17_Valid_Out, channel15_Kernel17_Valid_Out, channel16_Kernel17_Valid_Out, channel17_Kernel17_Valid_Out, channel18_Kernel17_Valid_Out, channel19_Kernel17_Valid_Out, channel20_Kernel17_Valid_Out, channel21_Kernel17_Valid_Out, channel22_Kernel17_Valid_Out, channel23_Kernel17_Valid_Out, channel24_Kernel17_Valid_Out, channel25_Kernel17_Valid_Out, channel26_Kernel17_Valid_Out, channel27_Kernel17_Valid_Out, channel28_Kernel17_Valid_Out, channel29_Kernel17_Valid_Out, channel30_Kernel17_Valid_Out, channel31_Kernel17_Valid_Out, channel32_Kernel17_Valid_Out;

	assign add_kernel17=channel1_Kernel17_Valid_Out & channel2_Kernel17_Valid_Out & channel3_Kernel17_Valid_Out & channel4_Kernel17_Valid_Out & channel5_Kernel17_Valid_Out & channel6_Kernel17_Valid_Out & channel7_Kernel17_Valid_Out & channel8_Kernel17_Valid_Out & channel9_Kernel17_Valid_Out & channel10_Kernel17_Valid_Out & channel11_Kernel17_Valid_Out & channel12_Kernel17_Valid_Out & channel13_Kernel17_Valid_Out & channel14_Kernel17_Valid_Out & channel15_Kernel17_Valid_Out & channel16_Kernel17_Valid_Out & channel17_Kernel17_Valid_Out & channel18_Kernel17_Valid_Out & channel19_Kernel17_Valid_Out & channel20_Kernel17_Valid_Out & channel21_Kernel17_Valid_Out & channel22_Kernel17_Valid_Out & channel23_Kernel17_Valid_Out & channel24_Kernel17_Valid_Out & channel25_Kernel17_Valid_Out & channel26_Kernel17_Valid_Out & channel27_Kernel17_Valid_Out & channel28_Kernel17_Valid_Out & channel29_Kernel17_Valid_Out & channel30_Kernel17_Valid_Out & channel31_Kernel17_Valid_Out & channel32_Kernel17_Valid_Out;

	wire channel1_Kernel18_Valid_Out, channel2_Kernel18_Valid_Out, channel3_Kernel18_Valid_Out, channel4_Kernel18_Valid_Out, channel5_Kernel18_Valid_Out, channel6_Kernel18_Valid_Out, channel7_Kernel18_Valid_Out, channel8_Kernel18_Valid_Out, channel9_Kernel18_Valid_Out, channel10_Kernel18_Valid_Out, channel11_Kernel18_Valid_Out, channel12_Kernel18_Valid_Out, channel13_Kernel18_Valid_Out, channel14_Kernel18_Valid_Out, channel15_Kernel18_Valid_Out, channel16_Kernel18_Valid_Out, channel17_Kernel18_Valid_Out, channel18_Kernel18_Valid_Out, channel19_Kernel18_Valid_Out, channel20_Kernel18_Valid_Out, channel21_Kernel18_Valid_Out, channel22_Kernel18_Valid_Out, channel23_Kernel18_Valid_Out, channel24_Kernel18_Valid_Out, channel25_Kernel18_Valid_Out, channel26_Kernel18_Valid_Out, channel27_Kernel18_Valid_Out, channel28_Kernel18_Valid_Out, channel29_Kernel18_Valid_Out, channel30_Kernel18_Valid_Out, channel31_Kernel18_Valid_Out, channel32_Kernel18_Valid_Out;

	assign add_kernel18=channel1_Kernel18_Valid_Out & channel2_Kernel18_Valid_Out & channel3_Kernel18_Valid_Out & channel4_Kernel18_Valid_Out & channel5_Kernel18_Valid_Out & channel6_Kernel18_Valid_Out & channel7_Kernel18_Valid_Out & channel8_Kernel18_Valid_Out & channel9_Kernel18_Valid_Out & channel10_Kernel18_Valid_Out & channel11_Kernel18_Valid_Out & channel12_Kernel18_Valid_Out & channel13_Kernel18_Valid_Out & channel14_Kernel18_Valid_Out & channel15_Kernel18_Valid_Out & channel16_Kernel18_Valid_Out & channel17_Kernel18_Valid_Out & channel18_Kernel18_Valid_Out & channel19_Kernel18_Valid_Out & channel20_Kernel18_Valid_Out & channel21_Kernel18_Valid_Out & channel22_Kernel18_Valid_Out & channel23_Kernel18_Valid_Out & channel24_Kernel18_Valid_Out & channel25_Kernel18_Valid_Out & channel26_Kernel18_Valid_Out & channel27_Kernel18_Valid_Out & channel28_Kernel18_Valid_Out & channel29_Kernel18_Valid_Out & channel30_Kernel18_Valid_Out & channel31_Kernel18_Valid_Out & channel32_Kernel18_Valid_Out;

	wire channel1_Kernel19_Valid_Out, channel2_Kernel19_Valid_Out, channel3_Kernel19_Valid_Out, channel4_Kernel19_Valid_Out, channel5_Kernel19_Valid_Out, channel6_Kernel19_Valid_Out, channel7_Kernel19_Valid_Out, channel8_Kernel19_Valid_Out, channel9_Kernel19_Valid_Out, channel10_Kernel19_Valid_Out, channel11_Kernel19_Valid_Out, channel12_Kernel19_Valid_Out, channel13_Kernel19_Valid_Out, channel14_Kernel19_Valid_Out, channel15_Kernel19_Valid_Out, channel16_Kernel19_Valid_Out, channel17_Kernel19_Valid_Out, channel18_Kernel19_Valid_Out, channel19_Kernel19_Valid_Out, channel20_Kernel19_Valid_Out, channel21_Kernel19_Valid_Out, channel22_Kernel19_Valid_Out, channel23_Kernel19_Valid_Out, channel24_Kernel19_Valid_Out, channel25_Kernel19_Valid_Out, channel26_Kernel19_Valid_Out, channel27_Kernel19_Valid_Out, channel28_Kernel19_Valid_Out, channel29_Kernel19_Valid_Out, channel30_Kernel19_Valid_Out, channel31_Kernel19_Valid_Out, channel32_Kernel19_Valid_Out;

	assign add_kernel19=channel1_Kernel19_Valid_Out & channel2_Kernel19_Valid_Out & channel3_Kernel19_Valid_Out & channel4_Kernel19_Valid_Out & channel5_Kernel19_Valid_Out & channel6_Kernel19_Valid_Out & channel7_Kernel19_Valid_Out & channel8_Kernel19_Valid_Out & channel9_Kernel19_Valid_Out & channel10_Kernel19_Valid_Out & channel11_Kernel19_Valid_Out & channel12_Kernel19_Valid_Out & channel13_Kernel19_Valid_Out & channel14_Kernel19_Valid_Out & channel15_Kernel19_Valid_Out & channel16_Kernel19_Valid_Out & channel17_Kernel19_Valid_Out & channel18_Kernel19_Valid_Out & channel19_Kernel19_Valid_Out & channel20_Kernel19_Valid_Out & channel21_Kernel19_Valid_Out & channel22_Kernel19_Valid_Out & channel23_Kernel19_Valid_Out & channel24_Kernel19_Valid_Out & channel25_Kernel19_Valid_Out & channel26_Kernel19_Valid_Out & channel27_Kernel19_Valid_Out & channel28_Kernel19_Valid_Out & channel29_Kernel19_Valid_Out & channel30_Kernel19_Valid_Out & channel31_Kernel19_Valid_Out & channel32_Kernel19_Valid_Out;

	wire channel1_Kernel20_Valid_Out, channel2_Kernel20_Valid_Out, channel3_Kernel20_Valid_Out, channel4_Kernel20_Valid_Out, channel5_Kernel20_Valid_Out, channel6_Kernel20_Valid_Out, channel7_Kernel20_Valid_Out, channel8_Kernel20_Valid_Out, channel9_Kernel20_Valid_Out, channel10_Kernel20_Valid_Out, channel11_Kernel20_Valid_Out, channel12_Kernel20_Valid_Out, channel13_Kernel20_Valid_Out, channel14_Kernel20_Valid_Out, channel15_Kernel20_Valid_Out, channel16_Kernel20_Valid_Out, channel17_Kernel20_Valid_Out, channel18_Kernel20_Valid_Out, channel19_Kernel20_Valid_Out, channel20_Kernel20_Valid_Out, channel21_Kernel20_Valid_Out, channel22_Kernel20_Valid_Out, channel23_Kernel20_Valid_Out, channel24_Kernel20_Valid_Out, channel25_Kernel20_Valid_Out, channel26_Kernel20_Valid_Out, channel27_Kernel20_Valid_Out, channel28_Kernel20_Valid_Out, channel29_Kernel20_Valid_Out, channel30_Kernel20_Valid_Out, channel31_Kernel20_Valid_Out, channel32_Kernel20_Valid_Out;

	assign add_kernel20=channel1_Kernel20_Valid_Out & channel2_Kernel20_Valid_Out & channel3_Kernel20_Valid_Out & channel4_Kernel20_Valid_Out & channel5_Kernel20_Valid_Out & channel6_Kernel20_Valid_Out & channel7_Kernel20_Valid_Out & channel8_Kernel20_Valid_Out & channel9_Kernel20_Valid_Out & channel10_Kernel20_Valid_Out & channel11_Kernel20_Valid_Out & channel12_Kernel20_Valid_Out & channel13_Kernel20_Valid_Out & channel14_Kernel20_Valid_Out & channel15_Kernel20_Valid_Out & channel16_Kernel20_Valid_Out & channel17_Kernel20_Valid_Out & channel18_Kernel20_Valid_Out & channel19_Kernel20_Valid_Out & channel20_Kernel20_Valid_Out & channel21_Kernel20_Valid_Out & channel22_Kernel20_Valid_Out & channel23_Kernel20_Valid_Out & channel24_Kernel20_Valid_Out & channel25_Kernel20_Valid_Out & channel26_Kernel20_Valid_Out & channel27_Kernel20_Valid_Out & channel28_Kernel20_Valid_Out & channel29_Kernel20_Valid_Out & channel30_Kernel20_Valid_Out & channel31_Kernel20_Valid_Out & channel32_Kernel20_Valid_Out;

	wire channel1_Kernel21_Valid_Out, channel2_Kernel21_Valid_Out, channel3_Kernel21_Valid_Out, channel4_Kernel21_Valid_Out, channel5_Kernel21_Valid_Out, channel6_Kernel21_Valid_Out, channel7_Kernel21_Valid_Out, channel8_Kernel21_Valid_Out, channel9_Kernel21_Valid_Out, channel10_Kernel21_Valid_Out, channel11_Kernel21_Valid_Out, channel12_Kernel21_Valid_Out, channel13_Kernel21_Valid_Out, channel14_Kernel21_Valid_Out, channel15_Kernel21_Valid_Out, channel16_Kernel21_Valid_Out, channel17_Kernel21_Valid_Out, channel18_Kernel21_Valid_Out, channel19_Kernel21_Valid_Out, channel20_Kernel21_Valid_Out, channel21_Kernel21_Valid_Out, channel22_Kernel21_Valid_Out, channel23_Kernel21_Valid_Out, channel24_Kernel21_Valid_Out, channel25_Kernel21_Valid_Out, channel26_Kernel21_Valid_Out, channel27_Kernel21_Valid_Out, channel28_Kernel21_Valid_Out, channel29_Kernel21_Valid_Out, channel30_Kernel21_Valid_Out, channel31_Kernel21_Valid_Out, channel32_Kernel21_Valid_Out;

	assign add_kernel21=channel1_Kernel21_Valid_Out & channel2_Kernel21_Valid_Out & channel3_Kernel21_Valid_Out & channel4_Kernel21_Valid_Out & channel5_Kernel21_Valid_Out & channel6_Kernel21_Valid_Out & channel7_Kernel21_Valid_Out & channel8_Kernel21_Valid_Out & channel9_Kernel21_Valid_Out & channel10_Kernel21_Valid_Out & channel11_Kernel21_Valid_Out & channel12_Kernel21_Valid_Out & channel13_Kernel21_Valid_Out & channel14_Kernel21_Valid_Out & channel15_Kernel21_Valid_Out & channel16_Kernel21_Valid_Out & channel17_Kernel21_Valid_Out & channel18_Kernel21_Valid_Out & channel19_Kernel21_Valid_Out & channel20_Kernel21_Valid_Out & channel21_Kernel21_Valid_Out & channel22_Kernel21_Valid_Out & channel23_Kernel21_Valid_Out & channel24_Kernel21_Valid_Out & channel25_Kernel21_Valid_Out & channel26_Kernel21_Valid_Out & channel27_Kernel21_Valid_Out & channel28_Kernel21_Valid_Out & channel29_Kernel21_Valid_Out & channel30_Kernel21_Valid_Out & channel31_Kernel21_Valid_Out & channel32_Kernel21_Valid_Out;

	wire channel1_Kernel22_Valid_Out, channel2_Kernel22_Valid_Out, channel3_Kernel22_Valid_Out, channel4_Kernel22_Valid_Out, channel5_Kernel22_Valid_Out, channel6_Kernel22_Valid_Out, channel7_Kernel22_Valid_Out, channel8_Kernel22_Valid_Out, channel9_Kernel22_Valid_Out, channel10_Kernel22_Valid_Out, channel11_Kernel22_Valid_Out, channel12_Kernel22_Valid_Out, channel13_Kernel22_Valid_Out, channel14_Kernel22_Valid_Out, channel15_Kernel22_Valid_Out, channel16_Kernel22_Valid_Out, channel17_Kernel22_Valid_Out, channel18_Kernel22_Valid_Out, channel19_Kernel22_Valid_Out, channel20_Kernel22_Valid_Out, channel21_Kernel22_Valid_Out, channel22_Kernel22_Valid_Out, channel23_Kernel22_Valid_Out, channel24_Kernel22_Valid_Out, channel25_Kernel22_Valid_Out, channel26_Kernel22_Valid_Out, channel27_Kernel22_Valid_Out, channel28_Kernel22_Valid_Out, channel29_Kernel22_Valid_Out, channel30_Kernel22_Valid_Out, channel31_Kernel22_Valid_Out, channel32_Kernel22_Valid_Out;

	assign add_kernel22=channel1_Kernel22_Valid_Out & channel2_Kernel22_Valid_Out & channel3_Kernel22_Valid_Out & channel4_Kernel22_Valid_Out & channel5_Kernel22_Valid_Out & channel6_Kernel22_Valid_Out & channel7_Kernel22_Valid_Out & channel8_Kernel22_Valid_Out & channel9_Kernel22_Valid_Out & channel10_Kernel22_Valid_Out & channel11_Kernel22_Valid_Out & channel12_Kernel22_Valid_Out & channel13_Kernel22_Valid_Out & channel14_Kernel22_Valid_Out & channel15_Kernel22_Valid_Out & channel16_Kernel22_Valid_Out & channel17_Kernel22_Valid_Out & channel18_Kernel22_Valid_Out & channel19_Kernel22_Valid_Out & channel20_Kernel22_Valid_Out & channel21_Kernel22_Valid_Out & channel22_Kernel22_Valid_Out & channel23_Kernel22_Valid_Out & channel24_Kernel22_Valid_Out & channel25_Kernel22_Valid_Out & channel26_Kernel22_Valid_Out & channel27_Kernel22_Valid_Out & channel28_Kernel22_Valid_Out & channel29_Kernel22_Valid_Out & channel30_Kernel22_Valid_Out & channel31_Kernel22_Valid_Out & channel32_Kernel22_Valid_Out;

	wire channel1_Kernel23_Valid_Out, channel2_Kernel23_Valid_Out, channel3_Kernel23_Valid_Out, channel4_Kernel23_Valid_Out, channel5_Kernel23_Valid_Out, channel6_Kernel23_Valid_Out, channel7_Kernel23_Valid_Out, channel8_Kernel23_Valid_Out, channel9_Kernel23_Valid_Out, channel10_Kernel23_Valid_Out, channel11_Kernel23_Valid_Out, channel12_Kernel23_Valid_Out, channel13_Kernel23_Valid_Out, channel14_Kernel23_Valid_Out, channel15_Kernel23_Valid_Out, channel16_Kernel23_Valid_Out, channel17_Kernel23_Valid_Out, channel18_Kernel23_Valid_Out, channel19_Kernel23_Valid_Out, channel20_Kernel23_Valid_Out, channel21_Kernel23_Valid_Out, channel22_Kernel23_Valid_Out, channel23_Kernel23_Valid_Out, channel24_Kernel23_Valid_Out, channel25_Kernel23_Valid_Out, channel26_Kernel23_Valid_Out, channel27_Kernel23_Valid_Out, channel28_Kernel23_Valid_Out, channel29_Kernel23_Valid_Out, channel30_Kernel23_Valid_Out, channel31_Kernel23_Valid_Out, channel32_Kernel23_Valid_Out;

	assign add_kernel23=channel1_Kernel23_Valid_Out & channel2_Kernel23_Valid_Out & channel3_Kernel23_Valid_Out & channel4_Kernel23_Valid_Out & channel5_Kernel23_Valid_Out & channel6_Kernel23_Valid_Out & channel7_Kernel23_Valid_Out & channel8_Kernel23_Valid_Out & channel9_Kernel23_Valid_Out & channel10_Kernel23_Valid_Out & channel11_Kernel23_Valid_Out & channel12_Kernel23_Valid_Out & channel13_Kernel23_Valid_Out & channel14_Kernel23_Valid_Out & channel15_Kernel23_Valid_Out & channel16_Kernel23_Valid_Out & channel17_Kernel23_Valid_Out & channel18_Kernel23_Valid_Out & channel19_Kernel23_Valid_Out & channel20_Kernel23_Valid_Out & channel21_Kernel23_Valid_Out & channel22_Kernel23_Valid_Out & channel23_Kernel23_Valid_Out & channel24_Kernel23_Valid_Out & channel25_Kernel23_Valid_Out & channel26_Kernel23_Valid_Out & channel27_Kernel23_Valid_Out & channel28_Kernel23_Valid_Out & channel29_Kernel23_Valid_Out & channel30_Kernel23_Valid_Out & channel31_Kernel23_Valid_Out & channel32_Kernel23_Valid_Out;

	wire channel1_Kernel24_Valid_Out, channel2_Kernel24_Valid_Out, channel3_Kernel24_Valid_Out, channel4_Kernel24_Valid_Out, channel5_Kernel24_Valid_Out, channel6_Kernel24_Valid_Out, channel7_Kernel24_Valid_Out, channel8_Kernel24_Valid_Out, channel9_Kernel24_Valid_Out, channel10_Kernel24_Valid_Out, channel11_Kernel24_Valid_Out, channel12_Kernel24_Valid_Out, channel13_Kernel24_Valid_Out, channel14_Kernel24_Valid_Out, channel15_Kernel24_Valid_Out, channel16_Kernel24_Valid_Out, channel17_Kernel24_Valid_Out, channel18_Kernel24_Valid_Out, channel19_Kernel24_Valid_Out, channel20_Kernel24_Valid_Out, channel21_Kernel24_Valid_Out, channel22_Kernel24_Valid_Out, channel23_Kernel24_Valid_Out, channel24_Kernel24_Valid_Out, channel25_Kernel24_Valid_Out, channel26_Kernel24_Valid_Out, channel27_Kernel24_Valid_Out, channel28_Kernel24_Valid_Out, channel29_Kernel24_Valid_Out, channel30_Kernel24_Valid_Out, channel31_Kernel24_Valid_Out, channel32_Kernel24_Valid_Out;

	assign add_kernel24=channel1_Kernel24_Valid_Out & channel2_Kernel24_Valid_Out & channel3_Kernel24_Valid_Out & channel4_Kernel24_Valid_Out & channel5_Kernel24_Valid_Out & channel6_Kernel24_Valid_Out & channel7_Kernel24_Valid_Out & channel8_Kernel24_Valid_Out & channel9_Kernel24_Valid_Out & channel10_Kernel24_Valid_Out & channel11_Kernel24_Valid_Out & channel12_Kernel24_Valid_Out & channel13_Kernel24_Valid_Out & channel14_Kernel24_Valid_Out & channel15_Kernel24_Valid_Out & channel16_Kernel24_Valid_Out & channel17_Kernel24_Valid_Out & channel18_Kernel24_Valid_Out & channel19_Kernel24_Valid_Out & channel20_Kernel24_Valid_Out & channel21_Kernel24_Valid_Out & channel22_Kernel24_Valid_Out & channel23_Kernel24_Valid_Out & channel24_Kernel24_Valid_Out & channel25_Kernel24_Valid_Out & channel26_Kernel24_Valid_Out & channel27_Kernel24_Valid_Out & channel28_Kernel24_Valid_Out & channel29_Kernel24_Valid_Out & channel30_Kernel24_Valid_Out & channel31_Kernel24_Valid_Out & channel32_Kernel24_Valid_Out;

	wire channel1_Kernel25_Valid_Out, channel2_Kernel25_Valid_Out, channel3_Kernel25_Valid_Out, channel4_Kernel25_Valid_Out, channel5_Kernel25_Valid_Out, channel6_Kernel25_Valid_Out, channel7_Kernel25_Valid_Out, channel8_Kernel25_Valid_Out, channel9_Kernel25_Valid_Out, channel10_Kernel25_Valid_Out, channel11_Kernel25_Valid_Out, channel12_Kernel25_Valid_Out, channel13_Kernel25_Valid_Out, channel14_Kernel25_Valid_Out, channel15_Kernel25_Valid_Out, channel16_Kernel25_Valid_Out, channel17_Kernel25_Valid_Out, channel18_Kernel25_Valid_Out, channel19_Kernel25_Valid_Out, channel20_Kernel25_Valid_Out, channel21_Kernel25_Valid_Out, channel22_Kernel25_Valid_Out, channel23_Kernel25_Valid_Out, channel24_Kernel25_Valid_Out, channel25_Kernel25_Valid_Out, channel26_Kernel25_Valid_Out, channel27_Kernel25_Valid_Out, channel28_Kernel25_Valid_Out, channel29_Kernel25_Valid_Out, channel30_Kernel25_Valid_Out, channel31_Kernel25_Valid_Out, channel32_Kernel25_Valid_Out;

	assign add_kernel25=channel1_Kernel25_Valid_Out & channel2_Kernel25_Valid_Out & channel3_Kernel25_Valid_Out & channel4_Kernel25_Valid_Out & channel5_Kernel25_Valid_Out & channel6_Kernel25_Valid_Out & channel7_Kernel25_Valid_Out & channel8_Kernel25_Valid_Out & channel9_Kernel25_Valid_Out & channel10_Kernel25_Valid_Out & channel11_Kernel25_Valid_Out & channel12_Kernel25_Valid_Out & channel13_Kernel25_Valid_Out & channel14_Kernel25_Valid_Out & channel15_Kernel25_Valid_Out & channel16_Kernel25_Valid_Out & channel17_Kernel25_Valid_Out & channel18_Kernel25_Valid_Out & channel19_Kernel25_Valid_Out & channel20_Kernel25_Valid_Out & channel21_Kernel25_Valid_Out & channel22_Kernel25_Valid_Out & channel23_Kernel25_Valid_Out & channel24_Kernel25_Valid_Out & channel25_Kernel25_Valid_Out & channel26_Kernel25_Valid_Out & channel27_Kernel25_Valid_Out & channel28_Kernel25_Valid_Out & channel29_Kernel25_Valid_Out & channel30_Kernel25_Valid_Out & channel31_Kernel25_Valid_Out & channel32_Kernel25_Valid_Out;

	wire channel1_Kernel26_Valid_Out, channel2_Kernel26_Valid_Out, channel3_Kernel26_Valid_Out, channel4_Kernel26_Valid_Out, channel5_Kernel26_Valid_Out, channel6_Kernel26_Valid_Out, channel7_Kernel26_Valid_Out, channel8_Kernel26_Valid_Out, channel9_Kernel26_Valid_Out, channel10_Kernel26_Valid_Out, channel11_Kernel26_Valid_Out, channel12_Kernel26_Valid_Out, channel13_Kernel26_Valid_Out, channel14_Kernel26_Valid_Out, channel15_Kernel26_Valid_Out, channel16_Kernel26_Valid_Out, channel17_Kernel26_Valid_Out, channel18_Kernel26_Valid_Out, channel19_Kernel26_Valid_Out, channel20_Kernel26_Valid_Out, channel21_Kernel26_Valid_Out, channel22_Kernel26_Valid_Out, channel23_Kernel26_Valid_Out, channel24_Kernel26_Valid_Out, channel25_Kernel26_Valid_Out, channel26_Kernel26_Valid_Out, channel27_Kernel26_Valid_Out, channel28_Kernel26_Valid_Out, channel29_Kernel26_Valid_Out, channel30_Kernel26_Valid_Out, channel31_Kernel26_Valid_Out, channel32_Kernel26_Valid_Out;

	assign add_kernel26=channel1_Kernel26_Valid_Out & channel2_Kernel26_Valid_Out & channel3_Kernel26_Valid_Out & channel4_Kernel26_Valid_Out & channel5_Kernel26_Valid_Out & channel6_Kernel26_Valid_Out & channel7_Kernel26_Valid_Out & channel8_Kernel26_Valid_Out & channel9_Kernel26_Valid_Out & channel10_Kernel26_Valid_Out & channel11_Kernel26_Valid_Out & channel12_Kernel26_Valid_Out & channel13_Kernel26_Valid_Out & channel14_Kernel26_Valid_Out & channel15_Kernel26_Valid_Out & channel16_Kernel26_Valid_Out & channel17_Kernel26_Valid_Out & channel18_Kernel26_Valid_Out & channel19_Kernel26_Valid_Out & channel20_Kernel26_Valid_Out & channel21_Kernel26_Valid_Out & channel22_Kernel26_Valid_Out & channel23_Kernel26_Valid_Out & channel24_Kernel26_Valid_Out & channel25_Kernel26_Valid_Out & channel26_Kernel26_Valid_Out & channel27_Kernel26_Valid_Out & channel28_Kernel26_Valid_Out & channel29_Kernel26_Valid_Out & channel30_Kernel26_Valid_Out & channel31_Kernel26_Valid_Out & channel32_Kernel26_Valid_Out;

	wire channel1_Kernel27_Valid_Out, channel2_Kernel27_Valid_Out, channel3_Kernel27_Valid_Out, channel4_Kernel27_Valid_Out, channel5_Kernel27_Valid_Out, channel6_Kernel27_Valid_Out, channel7_Kernel27_Valid_Out, channel8_Kernel27_Valid_Out, channel9_Kernel27_Valid_Out, channel10_Kernel27_Valid_Out, channel11_Kernel27_Valid_Out, channel12_Kernel27_Valid_Out, channel13_Kernel27_Valid_Out, channel14_Kernel27_Valid_Out, channel15_Kernel27_Valid_Out, channel16_Kernel27_Valid_Out, channel17_Kernel27_Valid_Out, channel18_Kernel27_Valid_Out, channel19_Kernel27_Valid_Out, channel20_Kernel27_Valid_Out, channel21_Kernel27_Valid_Out, channel22_Kernel27_Valid_Out, channel23_Kernel27_Valid_Out, channel24_Kernel27_Valid_Out, channel25_Kernel27_Valid_Out, channel26_Kernel27_Valid_Out, channel27_Kernel27_Valid_Out, channel28_Kernel27_Valid_Out, channel29_Kernel27_Valid_Out, channel30_Kernel27_Valid_Out, channel31_Kernel27_Valid_Out, channel32_Kernel27_Valid_Out;

	assign add_kernel27=channel1_Kernel27_Valid_Out & channel2_Kernel27_Valid_Out & channel3_Kernel27_Valid_Out & channel4_Kernel27_Valid_Out & channel5_Kernel27_Valid_Out & channel6_Kernel27_Valid_Out & channel7_Kernel27_Valid_Out & channel8_Kernel27_Valid_Out & channel9_Kernel27_Valid_Out & channel10_Kernel27_Valid_Out & channel11_Kernel27_Valid_Out & channel12_Kernel27_Valid_Out & channel13_Kernel27_Valid_Out & channel14_Kernel27_Valid_Out & channel15_Kernel27_Valid_Out & channel16_Kernel27_Valid_Out & channel17_Kernel27_Valid_Out & channel18_Kernel27_Valid_Out & channel19_Kernel27_Valid_Out & channel20_Kernel27_Valid_Out & channel21_Kernel27_Valid_Out & channel22_Kernel27_Valid_Out & channel23_Kernel27_Valid_Out & channel24_Kernel27_Valid_Out & channel25_Kernel27_Valid_Out & channel26_Kernel27_Valid_Out & channel27_Kernel27_Valid_Out & channel28_Kernel27_Valid_Out & channel29_Kernel27_Valid_Out & channel30_Kernel27_Valid_Out & channel31_Kernel27_Valid_Out & channel32_Kernel27_Valid_Out;

	wire channel1_Kernel28_Valid_Out, channel2_Kernel28_Valid_Out, channel3_Kernel28_Valid_Out, channel4_Kernel28_Valid_Out, channel5_Kernel28_Valid_Out, channel6_Kernel28_Valid_Out, channel7_Kernel28_Valid_Out, channel8_Kernel28_Valid_Out, channel9_Kernel28_Valid_Out, channel10_Kernel28_Valid_Out, channel11_Kernel28_Valid_Out, channel12_Kernel28_Valid_Out, channel13_Kernel28_Valid_Out, channel14_Kernel28_Valid_Out, channel15_Kernel28_Valid_Out, channel16_Kernel28_Valid_Out, channel17_Kernel28_Valid_Out, channel18_Kernel28_Valid_Out, channel19_Kernel28_Valid_Out, channel20_Kernel28_Valid_Out, channel21_Kernel28_Valid_Out, channel22_Kernel28_Valid_Out, channel23_Kernel28_Valid_Out, channel24_Kernel28_Valid_Out, channel25_Kernel28_Valid_Out, channel26_Kernel28_Valid_Out, channel27_Kernel28_Valid_Out, channel28_Kernel28_Valid_Out, channel29_Kernel28_Valid_Out, channel30_Kernel28_Valid_Out, channel31_Kernel28_Valid_Out, channel32_Kernel28_Valid_Out;

	assign add_kernel28=channel1_Kernel28_Valid_Out & channel2_Kernel28_Valid_Out & channel3_Kernel28_Valid_Out & channel4_Kernel28_Valid_Out & channel5_Kernel28_Valid_Out & channel6_Kernel28_Valid_Out & channel7_Kernel28_Valid_Out & channel8_Kernel28_Valid_Out & channel9_Kernel28_Valid_Out & channel10_Kernel28_Valid_Out & channel11_Kernel28_Valid_Out & channel12_Kernel28_Valid_Out & channel13_Kernel28_Valid_Out & channel14_Kernel28_Valid_Out & channel15_Kernel28_Valid_Out & channel16_Kernel28_Valid_Out & channel17_Kernel28_Valid_Out & channel18_Kernel28_Valid_Out & channel19_Kernel28_Valid_Out & channel20_Kernel28_Valid_Out & channel21_Kernel28_Valid_Out & channel22_Kernel28_Valid_Out & channel23_Kernel28_Valid_Out & channel24_Kernel28_Valid_Out & channel25_Kernel28_Valid_Out & channel26_Kernel28_Valid_Out & channel27_Kernel28_Valid_Out & channel28_Kernel28_Valid_Out & channel29_Kernel28_Valid_Out & channel30_Kernel28_Valid_Out & channel31_Kernel28_Valid_Out & channel32_Kernel28_Valid_Out;

	wire channel1_Kernel29_Valid_Out, channel2_Kernel29_Valid_Out, channel3_Kernel29_Valid_Out, channel4_Kernel29_Valid_Out, channel5_Kernel29_Valid_Out, channel6_Kernel29_Valid_Out, channel7_Kernel29_Valid_Out, channel8_Kernel29_Valid_Out, channel9_Kernel29_Valid_Out, channel10_Kernel29_Valid_Out, channel11_Kernel29_Valid_Out, channel12_Kernel29_Valid_Out, channel13_Kernel29_Valid_Out, channel14_Kernel29_Valid_Out, channel15_Kernel29_Valid_Out, channel16_Kernel29_Valid_Out, channel17_Kernel29_Valid_Out, channel18_Kernel29_Valid_Out, channel19_Kernel29_Valid_Out, channel20_Kernel29_Valid_Out, channel21_Kernel29_Valid_Out, channel22_Kernel29_Valid_Out, channel23_Kernel29_Valid_Out, channel24_Kernel29_Valid_Out, channel25_Kernel29_Valid_Out, channel26_Kernel29_Valid_Out, channel27_Kernel29_Valid_Out, channel28_Kernel29_Valid_Out, channel29_Kernel29_Valid_Out, channel30_Kernel29_Valid_Out, channel31_Kernel29_Valid_Out, channel32_Kernel29_Valid_Out;

	assign add_kernel29=channel1_Kernel29_Valid_Out & channel2_Kernel29_Valid_Out & channel3_Kernel29_Valid_Out & channel4_Kernel29_Valid_Out & channel5_Kernel29_Valid_Out & channel6_Kernel29_Valid_Out & channel7_Kernel29_Valid_Out & channel8_Kernel29_Valid_Out & channel9_Kernel29_Valid_Out & channel10_Kernel29_Valid_Out & channel11_Kernel29_Valid_Out & channel12_Kernel29_Valid_Out & channel13_Kernel29_Valid_Out & channel14_Kernel29_Valid_Out & channel15_Kernel29_Valid_Out & channel16_Kernel29_Valid_Out & channel17_Kernel29_Valid_Out & channel18_Kernel29_Valid_Out & channel19_Kernel29_Valid_Out & channel20_Kernel29_Valid_Out & channel21_Kernel29_Valid_Out & channel22_Kernel29_Valid_Out & channel23_Kernel29_Valid_Out & channel24_Kernel29_Valid_Out & channel25_Kernel29_Valid_Out & channel26_Kernel29_Valid_Out & channel27_Kernel29_Valid_Out & channel28_Kernel29_Valid_Out & channel29_Kernel29_Valid_Out & channel30_Kernel29_Valid_Out & channel31_Kernel29_Valid_Out & channel32_Kernel29_Valid_Out;

	wire channel1_Kernel30_Valid_Out, channel2_Kernel30_Valid_Out, channel3_Kernel30_Valid_Out, channel4_Kernel30_Valid_Out, channel5_Kernel30_Valid_Out, channel6_Kernel30_Valid_Out, channel7_Kernel30_Valid_Out, channel8_Kernel30_Valid_Out, channel9_Kernel30_Valid_Out, channel10_Kernel30_Valid_Out, channel11_Kernel30_Valid_Out, channel12_Kernel30_Valid_Out, channel13_Kernel30_Valid_Out, channel14_Kernel30_Valid_Out, channel15_Kernel30_Valid_Out, channel16_Kernel30_Valid_Out, channel17_Kernel30_Valid_Out, channel18_Kernel30_Valid_Out, channel19_Kernel30_Valid_Out, channel20_Kernel30_Valid_Out, channel21_Kernel30_Valid_Out, channel22_Kernel30_Valid_Out, channel23_Kernel30_Valid_Out, channel24_Kernel30_Valid_Out, channel25_Kernel30_Valid_Out, channel26_Kernel30_Valid_Out, channel27_Kernel30_Valid_Out, channel28_Kernel30_Valid_Out, channel29_Kernel30_Valid_Out, channel30_Kernel30_Valid_Out, channel31_Kernel30_Valid_Out, channel32_Kernel30_Valid_Out;

	assign add_kernel30=channel1_Kernel30_Valid_Out & channel2_Kernel30_Valid_Out & channel3_Kernel30_Valid_Out & channel4_Kernel30_Valid_Out & channel5_Kernel30_Valid_Out & channel6_Kernel30_Valid_Out & channel7_Kernel30_Valid_Out & channel8_Kernel30_Valid_Out & channel9_Kernel30_Valid_Out & channel10_Kernel30_Valid_Out & channel11_Kernel30_Valid_Out & channel12_Kernel30_Valid_Out & channel13_Kernel30_Valid_Out & channel14_Kernel30_Valid_Out & channel15_Kernel30_Valid_Out & channel16_Kernel30_Valid_Out & channel17_Kernel30_Valid_Out & channel18_Kernel30_Valid_Out & channel19_Kernel30_Valid_Out & channel20_Kernel30_Valid_Out & channel21_Kernel30_Valid_Out & channel22_Kernel30_Valid_Out & channel23_Kernel30_Valid_Out & channel24_Kernel30_Valid_Out & channel25_Kernel30_Valid_Out & channel26_Kernel30_Valid_Out & channel27_Kernel30_Valid_Out & channel28_Kernel30_Valid_Out & channel29_Kernel30_Valid_Out & channel30_Kernel30_Valid_Out & channel31_Kernel30_Valid_Out & channel32_Kernel30_Valid_Out;

	wire channel1_Kernel31_Valid_Out, channel2_Kernel31_Valid_Out, channel3_Kernel31_Valid_Out, channel4_Kernel31_Valid_Out, channel5_Kernel31_Valid_Out, channel6_Kernel31_Valid_Out, channel7_Kernel31_Valid_Out, channel8_Kernel31_Valid_Out, channel9_Kernel31_Valid_Out, channel10_Kernel31_Valid_Out, channel11_Kernel31_Valid_Out, channel12_Kernel31_Valid_Out, channel13_Kernel31_Valid_Out, channel14_Kernel31_Valid_Out, channel15_Kernel31_Valid_Out, channel16_Kernel31_Valid_Out, channel17_Kernel31_Valid_Out, channel18_Kernel31_Valid_Out, channel19_Kernel31_Valid_Out, channel20_Kernel31_Valid_Out, channel21_Kernel31_Valid_Out, channel22_Kernel31_Valid_Out, channel23_Kernel31_Valid_Out, channel24_Kernel31_Valid_Out, channel25_Kernel31_Valid_Out, channel26_Kernel31_Valid_Out, channel27_Kernel31_Valid_Out, channel28_Kernel31_Valid_Out, channel29_Kernel31_Valid_Out, channel30_Kernel31_Valid_Out, channel31_Kernel31_Valid_Out, channel32_Kernel31_Valid_Out;

	assign add_kernel31=channel1_Kernel31_Valid_Out & channel2_Kernel31_Valid_Out & channel3_Kernel31_Valid_Out & channel4_Kernel31_Valid_Out & channel5_Kernel31_Valid_Out & channel6_Kernel31_Valid_Out & channel7_Kernel31_Valid_Out & channel8_Kernel31_Valid_Out & channel9_Kernel31_Valid_Out & channel10_Kernel31_Valid_Out & channel11_Kernel31_Valid_Out & channel12_Kernel31_Valid_Out & channel13_Kernel31_Valid_Out & channel14_Kernel31_Valid_Out & channel15_Kernel31_Valid_Out & channel16_Kernel31_Valid_Out & channel17_Kernel31_Valid_Out & channel18_Kernel31_Valid_Out & channel19_Kernel31_Valid_Out & channel20_Kernel31_Valid_Out & channel21_Kernel31_Valid_Out & channel22_Kernel31_Valid_Out & channel23_Kernel31_Valid_Out & channel24_Kernel31_Valid_Out & channel25_Kernel31_Valid_Out & channel26_Kernel31_Valid_Out & channel27_Kernel31_Valid_Out & channel28_Kernel31_Valid_Out & channel29_Kernel31_Valid_Out & channel30_Kernel31_Valid_Out & channel31_Kernel31_Valid_Out & channel32_Kernel31_Valid_Out;

	wire channel1_Kernel32_Valid_Out, channel2_Kernel32_Valid_Out, channel3_Kernel32_Valid_Out, channel4_Kernel32_Valid_Out, channel5_Kernel32_Valid_Out, channel6_Kernel32_Valid_Out, channel7_Kernel32_Valid_Out, channel8_Kernel32_Valid_Out, channel9_Kernel32_Valid_Out, channel10_Kernel32_Valid_Out, channel11_Kernel32_Valid_Out, channel12_Kernel32_Valid_Out, channel13_Kernel32_Valid_Out, channel14_Kernel32_Valid_Out, channel15_Kernel32_Valid_Out, channel16_Kernel32_Valid_Out, channel17_Kernel32_Valid_Out, channel18_Kernel32_Valid_Out, channel19_Kernel32_Valid_Out, channel20_Kernel32_Valid_Out, channel21_Kernel32_Valid_Out, channel22_Kernel32_Valid_Out, channel23_Kernel32_Valid_Out, channel24_Kernel32_Valid_Out, channel25_Kernel32_Valid_Out, channel26_Kernel32_Valid_Out, channel27_Kernel32_Valid_Out, channel28_Kernel32_Valid_Out, channel29_Kernel32_Valid_Out, channel30_Kernel32_Valid_Out, channel31_Kernel32_Valid_Out, channel32_Kernel32_Valid_Out;

	assign add_kernel32=channel1_Kernel32_Valid_Out & channel2_Kernel32_Valid_Out & channel3_Kernel32_Valid_Out & channel4_Kernel32_Valid_Out & channel5_Kernel32_Valid_Out & channel6_Kernel32_Valid_Out & channel7_Kernel32_Valid_Out & channel8_Kernel32_Valid_Out & channel9_Kernel32_Valid_Out & channel10_Kernel32_Valid_Out & channel11_Kernel32_Valid_Out & channel12_Kernel32_Valid_Out & channel13_Kernel32_Valid_Out & channel14_Kernel32_Valid_Out & channel15_Kernel32_Valid_Out & channel16_Kernel32_Valid_Out & channel17_Kernel32_Valid_Out & channel18_Kernel32_Valid_Out & channel19_Kernel32_Valid_Out & channel20_Kernel32_Valid_Out & channel21_Kernel32_Valid_Out & channel22_Kernel32_Valid_Out & channel23_Kernel32_Valid_Out & channel24_Kernel32_Valid_Out & channel25_Kernel32_Valid_Out & channel26_Kernel32_Valid_Out & channel27_Kernel32_Valid_Out & channel28_Kernel32_Valid_Out & channel29_Kernel32_Valid_Out & channel30_Kernel32_Valid_Out & channel31_Kernel32_Valid_Out & channel32_Kernel32_Valid_Out;

	wire channel1_Kernel33_Valid_Out, channel2_Kernel33_Valid_Out, channel3_Kernel33_Valid_Out, channel4_Kernel33_Valid_Out, channel5_Kernel33_Valid_Out, channel6_Kernel33_Valid_Out, channel7_Kernel33_Valid_Out, channel8_Kernel33_Valid_Out, channel9_Kernel33_Valid_Out, channel10_Kernel33_Valid_Out, channel11_Kernel33_Valid_Out, channel12_Kernel33_Valid_Out, channel13_Kernel33_Valid_Out, channel14_Kernel33_Valid_Out, channel15_Kernel33_Valid_Out, channel16_Kernel33_Valid_Out, channel17_Kernel33_Valid_Out, channel18_Kernel33_Valid_Out, channel19_Kernel33_Valid_Out, channel20_Kernel33_Valid_Out, channel21_Kernel33_Valid_Out, channel22_Kernel33_Valid_Out, channel23_Kernel33_Valid_Out, channel24_Kernel33_Valid_Out, channel25_Kernel33_Valid_Out, channel26_Kernel33_Valid_Out, channel27_Kernel33_Valid_Out, channel28_Kernel33_Valid_Out, channel29_Kernel33_Valid_Out, channel30_Kernel33_Valid_Out, channel31_Kernel33_Valid_Out, channel32_Kernel33_Valid_Out;

	assign add_kernel33=channel1_Kernel33_Valid_Out & channel2_Kernel33_Valid_Out & channel3_Kernel33_Valid_Out & channel4_Kernel33_Valid_Out & channel5_Kernel33_Valid_Out & channel6_Kernel33_Valid_Out & channel7_Kernel33_Valid_Out & channel8_Kernel33_Valid_Out & channel9_Kernel33_Valid_Out & channel10_Kernel33_Valid_Out & channel11_Kernel33_Valid_Out & channel12_Kernel33_Valid_Out & channel13_Kernel33_Valid_Out & channel14_Kernel33_Valid_Out & channel15_Kernel33_Valid_Out & channel16_Kernel33_Valid_Out & channel17_Kernel33_Valid_Out & channel18_Kernel33_Valid_Out & channel19_Kernel33_Valid_Out & channel20_Kernel33_Valid_Out & channel21_Kernel33_Valid_Out & channel22_Kernel33_Valid_Out & channel23_Kernel33_Valid_Out & channel24_Kernel33_Valid_Out & channel25_Kernel33_Valid_Out & channel26_Kernel33_Valid_Out & channel27_Kernel33_Valid_Out & channel28_Kernel33_Valid_Out & channel29_Kernel33_Valid_Out & channel30_Kernel33_Valid_Out & channel31_Kernel33_Valid_Out & channel32_Kernel33_Valid_Out;

	wire channel1_Kernel34_Valid_Out, channel2_Kernel34_Valid_Out, channel3_Kernel34_Valid_Out, channel4_Kernel34_Valid_Out, channel5_Kernel34_Valid_Out, channel6_Kernel34_Valid_Out, channel7_Kernel34_Valid_Out, channel8_Kernel34_Valid_Out, channel9_Kernel34_Valid_Out, channel10_Kernel34_Valid_Out, channel11_Kernel34_Valid_Out, channel12_Kernel34_Valid_Out, channel13_Kernel34_Valid_Out, channel14_Kernel34_Valid_Out, channel15_Kernel34_Valid_Out, channel16_Kernel34_Valid_Out, channel17_Kernel34_Valid_Out, channel18_Kernel34_Valid_Out, channel19_Kernel34_Valid_Out, channel20_Kernel34_Valid_Out, channel21_Kernel34_Valid_Out, channel22_Kernel34_Valid_Out, channel23_Kernel34_Valid_Out, channel24_Kernel34_Valid_Out, channel25_Kernel34_Valid_Out, channel26_Kernel34_Valid_Out, channel27_Kernel34_Valid_Out, channel28_Kernel34_Valid_Out, channel29_Kernel34_Valid_Out, channel30_Kernel34_Valid_Out, channel31_Kernel34_Valid_Out, channel32_Kernel34_Valid_Out;

	assign add_kernel34=channel1_Kernel34_Valid_Out & channel2_Kernel34_Valid_Out & channel3_Kernel34_Valid_Out & channel4_Kernel34_Valid_Out & channel5_Kernel34_Valid_Out & channel6_Kernel34_Valid_Out & channel7_Kernel34_Valid_Out & channel8_Kernel34_Valid_Out & channel9_Kernel34_Valid_Out & channel10_Kernel34_Valid_Out & channel11_Kernel34_Valid_Out & channel12_Kernel34_Valid_Out & channel13_Kernel34_Valid_Out & channel14_Kernel34_Valid_Out & channel15_Kernel34_Valid_Out & channel16_Kernel34_Valid_Out & channel17_Kernel34_Valid_Out & channel18_Kernel34_Valid_Out & channel19_Kernel34_Valid_Out & channel20_Kernel34_Valid_Out & channel21_Kernel34_Valid_Out & channel22_Kernel34_Valid_Out & channel23_Kernel34_Valid_Out & channel24_Kernel34_Valid_Out & channel25_Kernel34_Valid_Out & channel26_Kernel34_Valid_Out & channel27_Kernel34_Valid_Out & channel28_Kernel34_Valid_Out & channel29_Kernel34_Valid_Out & channel30_Kernel34_Valid_Out & channel31_Kernel34_Valid_Out & channel32_Kernel34_Valid_Out;

	wire channel1_Kernel35_Valid_Out, channel2_Kernel35_Valid_Out, channel3_Kernel35_Valid_Out, channel4_Kernel35_Valid_Out, channel5_Kernel35_Valid_Out, channel6_Kernel35_Valid_Out, channel7_Kernel35_Valid_Out, channel8_Kernel35_Valid_Out, channel9_Kernel35_Valid_Out, channel10_Kernel35_Valid_Out, channel11_Kernel35_Valid_Out, channel12_Kernel35_Valid_Out, channel13_Kernel35_Valid_Out, channel14_Kernel35_Valid_Out, channel15_Kernel35_Valid_Out, channel16_Kernel35_Valid_Out, channel17_Kernel35_Valid_Out, channel18_Kernel35_Valid_Out, channel19_Kernel35_Valid_Out, channel20_Kernel35_Valid_Out, channel21_Kernel35_Valid_Out, channel22_Kernel35_Valid_Out, channel23_Kernel35_Valid_Out, channel24_Kernel35_Valid_Out, channel25_Kernel35_Valid_Out, channel26_Kernel35_Valid_Out, channel27_Kernel35_Valid_Out, channel28_Kernel35_Valid_Out, channel29_Kernel35_Valid_Out, channel30_Kernel35_Valid_Out, channel31_Kernel35_Valid_Out, channel32_Kernel35_Valid_Out;

	assign add_kernel35=channel1_Kernel35_Valid_Out & channel2_Kernel35_Valid_Out & channel3_Kernel35_Valid_Out & channel4_Kernel35_Valid_Out & channel5_Kernel35_Valid_Out & channel6_Kernel35_Valid_Out & channel7_Kernel35_Valid_Out & channel8_Kernel35_Valid_Out & channel9_Kernel35_Valid_Out & channel10_Kernel35_Valid_Out & channel11_Kernel35_Valid_Out & channel12_Kernel35_Valid_Out & channel13_Kernel35_Valid_Out & channel14_Kernel35_Valid_Out & channel15_Kernel35_Valid_Out & channel16_Kernel35_Valid_Out & channel17_Kernel35_Valid_Out & channel18_Kernel35_Valid_Out & channel19_Kernel35_Valid_Out & channel20_Kernel35_Valid_Out & channel21_Kernel35_Valid_Out & channel22_Kernel35_Valid_Out & channel23_Kernel35_Valid_Out & channel24_Kernel35_Valid_Out & channel25_Kernel35_Valid_Out & channel26_Kernel35_Valid_Out & channel27_Kernel35_Valid_Out & channel28_Kernel35_Valid_Out & channel29_Kernel35_Valid_Out & channel30_Kernel35_Valid_Out & channel31_Kernel35_Valid_Out & channel32_Kernel35_Valid_Out;

	wire channel1_Kernel36_Valid_Out, channel2_Kernel36_Valid_Out, channel3_Kernel36_Valid_Out, channel4_Kernel36_Valid_Out, channel5_Kernel36_Valid_Out, channel6_Kernel36_Valid_Out, channel7_Kernel36_Valid_Out, channel8_Kernel36_Valid_Out, channel9_Kernel36_Valid_Out, channel10_Kernel36_Valid_Out, channel11_Kernel36_Valid_Out, channel12_Kernel36_Valid_Out, channel13_Kernel36_Valid_Out, channel14_Kernel36_Valid_Out, channel15_Kernel36_Valid_Out, channel16_Kernel36_Valid_Out, channel17_Kernel36_Valid_Out, channel18_Kernel36_Valid_Out, channel19_Kernel36_Valid_Out, channel20_Kernel36_Valid_Out, channel21_Kernel36_Valid_Out, channel22_Kernel36_Valid_Out, channel23_Kernel36_Valid_Out, channel24_Kernel36_Valid_Out, channel25_Kernel36_Valid_Out, channel26_Kernel36_Valid_Out, channel27_Kernel36_Valid_Out, channel28_Kernel36_Valid_Out, channel29_Kernel36_Valid_Out, channel30_Kernel36_Valid_Out, channel31_Kernel36_Valid_Out, channel32_Kernel36_Valid_Out;

	assign add_kernel36=channel1_Kernel36_Valid_Out & channel2_Kernel36_Valid_Out & channel3_Kernel36_Valid_Out & channel4_Kernel36_Valid_Out & channel5_Kernel36_Valid_Out & channel6_Kernel36_Valid_Out & channel7_Kernel36_Valid_Out & channel8_Kernel36_Valid_Out & channel9_Kernel36_Valid_Out & channel10_Kernel36_Valid_Out & channel11_Kernel36_Valid_Out & channel12_Kernel36_Valid_Out & channel13_Kernel36_Valid_Out & channel14_Kernel36_Valid_Out & channel15_Kernel36_Valid_Out & channel16_Kernel36_Valid_Out & channel17_Kernel36_Valid_Out & channel18_Kernel36_Valid_Out & channel19_Kernel36_Valid_Out & channel20_Kernel36_Valid_Out & channel21_Kernel36_Valid_Out & channel22_Kernel36_Valid_Out & channel23_Kernel36_Valid_Out & channel24_Kernel36_Valid_Out & channel25_Kernel36_Valid_Out & channel26_Kernel36_Valid_Out & channel27_Kernel36_Valid_Out & channel28_Kernel36_Valid_Out & channel29_Kernel36_Valid_Out & channel30_Kernel36_Valid_Out & channel31_Kernel36_Valid_Out & channel32_Kernel36_Valid_Out;

	wire channel1_Kernel37_Valid_Out, channel2_Kernel37_Valid_Out, channel3_Kernel37_Valid_Out, channel4_Kernel37_Valid_Out, channel5_Kernel37_Valid_Out, channel6_Kernel37_Valid_Out, channel7_Kernel37_Valid_Out, channel8_Kernel37_Valid_Out, channel9_Kernel37_Valid_Out, channel10_Kernel37_Valid_Out, channel11_Kernel37_Valid_Out, channel12_Kernel37_Valid_Out, channel13_Kernel37_Valid_Out, channel14_Kernel37_Valid_Out, channel15_Kernel37_Valid_Out, channel16_Kernel37_Valid_Out, channel17_Kernel37_Valid_Out, channel18_Kernel37_Valid_Out, channel19_Kernel37_Valid_Out, channel20_Kernel37_Valid_Out, channel21_Kernel37_Valid_Out, channel22_Kernel37_Valid_Out, channel23_Kernel37_Valid_Out, channel24_Kernel37_Valid_Out, channel25_Kernel37_Valid_Out, channel26_Kernel37_Valid_Out, channel27_Kernel37_Valid_Out, channel28_Kernel37_Valid_Out, channel29_Kernel37_Valid_Out, channel30_Kernel37_Valid_Out, channel31_Kernel37_Valid_Out, channel32_Kernel37_Valid_Out;

	assign add_kernel37=channel1_Kernel37_Valid_Out & channel2_Kernel37_Valid_Out & channel3_Kernel37_Valid_Out & channel4_Kernel37_Valid_Out & channel5_Kernel37_Valid_Out & channel6_Kernel37_Valid_Out & channel7_Kernel37_Valid_Out & channel8_Kernel37_Valid_Out & channel9_Kernel37_Valid_Out & channel10_Kernel37_Valid_Out & channel11_Kernel37_Valid_Out & channel12_Kernel37_Valid_Out & channel13_Kernel37_Valid_Out & channel14_Kernel37_Valid_Out & channel15_Kernel37_Valid_Out & channel16_Kernel37_Valid_Out & channel17_Kernel37_Valid_Out & channel18_Kernel37_Valid_Out & channel19_Kernel37_Valid_Out & channel20_Kernel37_Valid_Out & channel21_Kernel37_Valid_Out & channel22_Kernel37_Valid_Out & channel23_Kernel37_Valid_Out & channel24_Kernel37_Valid_Out & channel25_Kernel37_Valid_Out & channel26_Kernel37_Valid_Out & channel27_Kernel37_Valid_Out & channel28_Kernel37_Valid_Out & channel29_Kernel37_Valid_Out & channel30_Kernel37_Valid_Out & channel31_Kernel37_Valid_Out & channel32_Kernel37_Valid_Out;

	wire channel1_Kernel38_Valid_Out, channel2_Kernel38_Valid_Out, channel3_Kernel38_Valid_Out, channel4_Kernel38_Valid_Out, channel5_Kernel38_Valid_Out, channel6_Kernel38_Valid_Out, channel7_Kernel38_Valid_Out, channel8_Kernel38_Valid_Out, channel9_Kernel38_Valid_Out, channel10_Kernel38_Valid_Out, channel11_Kernel38_Valid_Out, channel12_Kernel38_Valid_Out, channel13_Kernel38_Valid_Out, channel14_Kernel38_Valid_Out, channel15_Kernel38_Valid_Out, channel16_Kernel38_Valid_Out, channel17_Kernel38_Valid_Out, channel18_Kernel38_Valid_Out, channel19_Kernel38_Valid_Out, channel20_Kernel38_Valid_Out, channel21_Kernel38_Valid_Out, channel22_Kernel38_Valid_Out, channel23_Kernel38_Valid_Out, channel24_Kernel38_Valid_Out, channel25_Kernel38_Valid_Out, channel26_Kernel38_Valid_Out, channel27_Kernel38_Valid_Out, channel28_Kernel38_Valid_Out, channel29_Kernel38_Valid_Out, channel30_Kernel38_Valid_Out, channel31_Kernel38_Valid_Out, channel32_Kernel38_Valid_Out;

	assign add_kernel38=channel1_Kernel38_Valid_Out & channel2_Kernel38_Valid_Out & channel3_Kernel38_Valid_Out & channel4_Kernel38_Valid_Out & channel5_Kernel38_Valid_Out & channel6_Kernel38_Valid_Out & channel7_Kernel38_Valid_Out & channel8_Kernel38_Valid_Out & channel9_Kernel38_Valid_Out & channel10_Kernel38_Valid_Out & channel11_Kernel38_Valid_Out & channel12_Kernel38_Valid_Out & channel13_Kernel38_Valid_Out & channel14_Kernel38_Valid_Out & channel15_Kernel38_Valid_Out & channel16_Kernel38_Valid_Out & channel17_Kernel38_Valid_Out & channel18_Kernel38_Valid_Out & channel19_Kernel38_Valid_Out & channel20_Kernel38_Valid_Out & channel21_Kernel38_Valid_Out & channel22_Kernel38_Valid_Out & channel23_Kernel38_Valid_Out & channel24_Kernel38_Valid_Out & channel25_Kernel38_Valid_Out & channel26_Kernel38_Valid_Out & channel27_Kernel38_Valid_Out & channel28_Kernel38_Valid_Out & channel29_Kernel38_Valid_Out & channel30_Kernel38_Valid_Out & channel31_Kernel38_Valid_Out & channel32_Kernel38_Valid_Out;

	wire channel1_Kernel39_Valid_Out, channel2_Kernel39_Valid_Out, channel3_Kernel39_Valid_Out, channel4_Kernel39_Valid_Out, channel5_Kernel39_Valid_Out, channel6_Kernel39_Valid_Out, channel7_Kernel39_Valid_Out, channel8_Kernel39_Valid_Out, channel9_Kernel39_Valid_Out, channel10_Kernel39_Valid_Out, channel11_Kernel39_Valid_Out, channel12_Kernel39_Valid_Out, channel13_Kernel39_Valid_Out, channel14_Kernel39_Valid_Out, channel15_Kernel39_Valid_Out, channel16_Kernel39_Valid_Out, channel17_Kernel39_Valid_Out, channel18_Kernel39_Valid_Out, channel19_Kernel39_Valid_Out, channel20_Kernel39_Valid_Out, channel21_Kernel39_Valid_Out, channel22_Kernel39_Valid_Out, channel23_Kernel39_Valid_Out, channel24_Kernel39_Valid_Out, channel25_Kernel39_Valid_Out, channel26_Kernel39_Valid_Out, channel27_Kernel39_Valid_Out, channel28_Kernel39_Valid_Out, channel29_Kernel39_Valid_Out, channel30_Kernel39_Valid_Out, channel31_Kernel39_Valid_Out, channel32_Kernel39_Valid_Out;

	assign add_kernel39=channel1_Kernel39_Valid_Out & channel2_Kernel39_Valid_Out & channel3_Kernel39_Valid_Out & channel4_Kernel39_Valid_Out & channel5_Kernel39_Valid_Out & channel6_Kernel39_Valid_Out & channel7_Kernel39_Valid_Out & channel8_Kernel39_Valid_Out & channel9_Kernel39_Valid_Out & channel10_Kernel39_Valid_Out & channel11_Kernel39_Valid_Out & channel12_Kernel39_Valid_Out & channel13_Kernel39_Valid_Out & channel14_Kernel39_Valid_Out & channel15_Kernel39_Valid_Out & channel16_Kernel39_Valid_Out & channel17_Kernel39_Valid_Out & channel18_Kernel39_Valid_Out & channel19_Kernel39_Valid_Out & channel20_Kernel39_Valid_Out & channel21_Kernel39_Valid_Out & channel22_Kernel39_Valid_Out & channel23_Kernel39_Valid_Out & channel24_Kernel39_Valid_Out & channel25_Kernel39_Valid_Out & channel26_Kernel39_Valid_Out & channel27_Kernel39_Valid_Out & channel28_Kernel39_Valid_Out & channel29_Kernel39_Valid_Out & channel30_Kernel39_Valid_Out & channel31_Kernel39_Valid_Out & channel32_Kernel39_Valid_Out;

	wire channel1_Kernel40_Valid_Out, channel2_Kernel40_Valid_Out, channel3_Kernel40_Valid_Out, channel4_Kernel40_Valid_Out, channel5_Kernel40_Valid_Out, channel6_Kernel40_Valid_Out, channel7_Kernel40_Valid_Out, channel8_Kernel40_Valid_Out, channel9_Kernel40_Valid_Out, channel10_Kernel40_Valid_Out, channel11_Kernel40_Valid_Out, channel12_Kernel40_Valid_Out, channel13_Kernel40_Valid_Out, channel14_Kernel40_Valid_Out, channel15_Kernel40_Valid_Out, channel16_Kernel40_Valid_Out, channel17_Kernel40_Valid_Out, channel18_Kernel40_Valid_Out, channel19_Kernel40_Valid_Out, channel20_Kernel40_Valid_Out, channel21_Kernel40_Valid_Out, channel22_Kernel40_Valid_Out, channel23_Kernel40_Valid_Out, channel24_Kernel40_Valid_Out, channel25_Kernel40_Valid_Out, channel26_Kernel40_Valid_Out, channel27_Kernel40_Valid_Out, channel28_Kernel40_Valid_Out, channel29_Kernel40_Valid_Out, channel30_Kernel40_Valid_Out, channel31_Kernel40_Valid_Out, channel32_Kernel40_Valid_Out;

	assign add_kernel40=channel1_Kernel40_Valid_Out & channel2_Kernel40_Valid_Out & channel3_Kernel40_Valid_Out & channel4_Kernel40_Valid_Out & channel5_Kernel40_Valid_Out & channel6_Kernel40_Valid_Out & channel7_Kernel40_Valid_Out & channel8_Kernel40_Valid_Out & channel9_Kernel40_Valid_Out & channel10_Kernel40_Valid_Out & channel11_Kernel40_Valid_Out & channel12_Kernel40_Valid_Out & channel13_Kernel40_Valid_Out & channel14_Kernel40_Valid_Out & channel15_Kernel40_Valid_Out & channel16_Kernel40_Valid_Out & channel17_Kernel40_Valid_Out & channel18_Kernel40_Valid_Out & channel19_Kernel40_Valid_Out & channel20_Kernel40_Valid_Out & channel21_Kernel40_Valid_Out & channel22_Kernel40_Valid_Out & channel23_Kernel40_Valid_Out & channel24_Kernel40_Valid_Out & channel25_Kernel40_Valid_Out & channel26_Kernel40_Valid_Out & channel27_Kernel40_Valid_Out & channel28_Kernel40_Valid_Out & channel29_Kernel40_Valid_Out & channel30_Kernel40_Valid_Out & channel31_Kernel40_Valid_Out & channel32_Kernel40_Valid_Out;

	wire channel1_Kernel41_Valid_Out, channel2_Kernel41_Valid_Out, channel3_Kernel41_Valid_Out, channel4_Kernel41_Valid_Out, channel5_Kernel41_Valid_Out, channel6_Kernel41_Valid_Out, channel7_Kernel41_Valid_Out, channel8_Kernel41_Valid_Out, channel9_Kernel41_Valid_Out, channel10_Kernel41_Valid_Out, channel11_Kernel41_Valid_Out, channel12_Kernel41_Valid_Out, channel13_Kernel41_Valid_Out, channel14_Kernel41_Valid_Out, channel15_Kernel41_Valid_Out, channel16_Kernel41_Valid_Out, channel17_Kernel41_Valid_Out, channel18_Kernel41_Valid_Out, channel19_Kernel41_Valid_Out, channel20_Kernel41_Valid_Out, channel21_Kernel41_Valid_Out, channel22_Kernel41_Valid_Out, channel23_Kernel41_Valid_Out, channel24_Kernel41_Valid_Out, channel25_Kernel41_Valid_Out, channel26_Kernel41_Valid_Out, channel27_Kernel41_Valid_Out, channel28_Kernel41_Valid_Out, channel29_Kernel41_Valid_Out, channel30_Kernel41_Valid_Out, channel31_Kernel41_Valid_Out, channel32_Kernel41_Valid_Out;

	assign add_kernel41=channel1_Kernel41_Valid_Out & channel2_Kernel41_Valid_Out & channel3_Kernel41_Valid_Out & channel4_Kernel41_Valid_Out & channel5_Kernel41_Valid_Out & channel6_Kernel41_Valid_Out & channel7_Kernel41_Valid_Out & channel8_Kernel41_Valid_Out & channel9_Kernel41_Valid_Out & channel10_Kernel41_Valid_Out & channel11_Kernel41_Valid_Out & channel12_Kernel41_Valid_Out & channel13_Kernel41_Valid_Out & channel14_Kernel41_Valid_Out & channel15_Kernel41_Valid_Out & channel16_Kernel41_Valid_Out & channel17_Kernel41_Valid_Out & channel18_Kernel41_Valid_Out & channel19_Kernel41_Valid_Out & channel20_Kernel41_Valid_Out & channel21_Kernel41_Valid_Out & channel22_Kernel41_Valid_Out & channel23_Kernel41_Valid_Out & channel24_Kernel41_Valid_Out & channel25_Kernel41_Valid_Out & channel26_Kernel41_Valid_Out & channel27_Kernel41_Valid_Out & channel28_Kernel41_Valid_Out & channel29_Kernel41_Valid_Out & channel30_Kernel41_Valid_Out & channel31_Kernel41_Valid_Out & channel32_Kernel41_Valid_Out;

	wire channel1_Kernel42_Valid_Out, channel2_Kernel42_Valid_Out, channel3_Kernel42_Valid_Out, channel4_Kernel42_Valid_Out, channel5_Kernel42_Valid_Out, channel6_Kernel42_Valid_Out, channel7_Kernel42_Valid_Out, channel8_Kernel42_Valid_Out, channel9_Kernel42_Valid_Out, channel10_Kernel42_Valid_Out, channel11_Kernel42_Valid_Out, channel12_Kernel42_Valid_Out, channel13_Kernel42_Valid_Out, channel14_Kernel42_Valid_Out, channel15_Kernel42_Valid_Out, channel16_Kernel42_Valid_Out, channel17_Kernel42_Valid_Out, channel18_Kernel42_Valid_Out, channel19_Kernel42_Valid_Out, channel20_Kernel42_Valid_Out, channel21_Kernel42_Valid_Out, channel22_Kernel42_Valid_Out, channel23_Kernel42_Valid_Out, channel24_Kernel42_Valid_Out, channel25_Kernel42_Valid_Out, channel26_Kernel42_Valid_Out, channel27_Kernel42_Valid_Out, channel28_Kernel42_Valid_Out, channel29_Kernel42_Valid_Out, channel30_Kernel42_Valid_Out, channel31_Kernel42_Valid_Out, channel32_Kernel42_Valid_Out;

	assign add_kernel42=channel1_Kernel42_Valid_Out & channel2_Kernel42_Valid_Out & channel3_Kernel42_Valid_Out & channel4_Kernel42_Valid_Out & channel5_Kernel42_Valid_Out & channel6_Kernel42_Valid_Out & channel7_Kernel42_Valid_Out & channel8_Kernel42_Valid_Out & channel9_Kernel42_Valid_Out & channel10_Kernel42_Valid_Out & channel11_Kernel42_Valid_Out & channel12_Kernel42_Valid_Out & channel13_Kernel42_Valid_Out & channel14_Kernel42_Valid_Out & channel15_Kernel42_Valid_Out & channel16_Kernel42_Valid_Out & channel17_Kernel42_Valid_Out & channel18_Kernel42_Valid_Out & channel19_Kernel42_Valid_Out & channel20_Kernel42_Valid_Out & channel21_Kernel42_Valid_Out & channel22_Kernel42_Valid_Out & channel23_Kernel42_Valid_Out & channel24_Kernel42_Valid_Out & channel25_Kernel42_Valid_Out & channel26_Kernel42_Valid_Out & channel27_Kernel42_Valid_Out & channel28_Kernel42_Valid_Out & channel29_Kernel42_Valid_Out & channel30_Kernel42_Valid_Out & channel31_Kernel42_Valid_Out & channel32_Kernel42_Valid_Out;

	wire channel1_Kernel43_Valid_Out, channel2_Kernel43_Valid_Out, channel3_Kernel43_Valid_Out, channel4_Kernel43_Valid_Out, channel5_Kernel43_Valid_Out, channel6_Kernel43_Valid_Out, channel7_Kernel43_Valid_Out, channel8_Kernel43_Valid_Out, channel9_Kernel43_Valid_Out, channel10_Kernel43_Valid_Out, channel11_Kernel43_Valid_Out, channel12_Kernel43_Valid_Out, channel13_Kernel43_Valid_Out, channel14_Kernel43_Valid_Out, channel15_Kernel43_Valid_Out, channel16_Kernel43_Valid_Out, channel17_Kernel43_Valid_Out, channel18_Kernel43_Valid_Out, channel19_Kernel43_Valid_Out, channel20_Kernel43_Valid_Out, channel21_Kernel43_Valid_Out, channel22_Kernel43_Valid_Out, channel23_Kernel43_Valid_Out, channel24_Kernel43_Valid_Out, channel25_Kernel43_Valid_Out, channel26_Kernel43_Valid_Out, channel27_Kernel43_Valid_Out, channel28_Kernel43_Valid_Out, channel29_Kernel43_Valid_Out, channel30_Kernel43_Valid_Out, channel31_Kernel43_Valid_Out, channel32_Kernel43_Valid_Out;

	assign add_kernel43=channel1_Kernel43_Valid_Out & channel2_Kernel43_Valid_Out & channel3_Kernel43_Valid_Out & channel4_Kernel43_Valid_Out & channel5_Kernel43_Valid_Out & channel6_Kernel43_Valid_Out & channel7_Kernel43_Valid_Out & channel8_Kernel43_Valid_Out & channel9_Kernel43_Valid_Out & channel10_Kernel43_Valid_Out & channel11_Kernel43_Valid_Out & channel12_Kernel43_Valid_Out & channel13_Kernel43_Valid_Out & channel14_Kernel43_Valid_Out & channel15_Kernel43_Valid_Out & channel16_Kernel43_Valid_Out & channel17_Kernel43_Valid_Out & channel18_Kernel43_Valid_Out & channel19_Kernel43_Valid_Out & channel20_Kernel43_Valid_Out & channel21_Kernel43_Valid_Out & channel22_Kernel43_Valid_Out & channel23_Kernel43_Valid_Out & channel24_Kernel43_Valid_Out & channel25_Kernel43_Valid_Out & channel26_Kernel43_Valid_Out & channel27_Kernel43_Valid_Out & channel28_Kernel43_Valid_Out & channel29_Kernel43_Valid_Out & channel30_Kernel43_Valid_Out & channel31_Kernel43_Valid_Out & channel32_Kernel43_Valid_Out;

	wire channel1_Kernel44_Valid_Out, channel2_Kernel44_Valid_Out, channel3_Kernel44_Valid_Out, channel4_Kernel44_Valid_Out, channel5_Kernel44_Valid_Out, channel6_Kernel44_Valid_Out, channel7_Kernel44_Valid_Out, channel8_Kernel44_Valid_Out, channel9_Kernel44_Valid_Out, channel10_Kernel44_Valid_Out, channel11_Kernel44_Valid_Out, channel12_Kernel44_Valid_Out, channel13_Kernel44_Valid_Out, channel14_Kernel44_Valid_Out, channel15_Kernel44_Valid_Out, channel16_Kernel44_Valid_Out, channel17_Kernel44_Valid_Out, channel18_Kernel44_Valid_Out, channel19_Kernel44_Valid_Out, channel20_Kernel44_Valid_Out, channel21_Kernel44_Valid_Out, channel22_Kernel44_Valid_Out, channel23_Kernel44_Valid_Out, channel24_Kernel44_Valid_Out, channel25_Kernel44_Valid_Out, channel26_Kernel44_Valid_Out, channel27_Kernel44_Valid_Out, channel28_Kernel44_Valid_Out, channel29_Kernel44_Valid_Out, channel30_Kernel44_Valid_Out, channel31_Kernel44_Valid_Out, channel32_Kernel44_Valid_Out;

	assign add_kernel44=channel1_Kernel44_Valid_Out & channel2_Kernel44_Valid_Out & channel3_Kernel44_Valid_Out & channel4_Kernel44_Valid_Out & channel5_Kernel44_Valid_Out & channel6_Kernel44_Valid_Out & channel7_Kernel44_Valid_Out & channel8_Kernel44_Valid_Out & channel9_Kernel44_Valid_Out & channel10_Kernel44_Valid_Out & channel11_Kernel44_Valid_Out & channel12_Kernel44_Valid_Out & channel13_Kernel44_Valid_Out & channel14_Kernel44_Valid_Out & channel15_Kernel44_Valid_Out & channel16_Kernel44_Valid_Out & channel17_Kernel44_Valid_Out & channel18_Kernel44_Valid_Out & channel19_Kernel44_Valid_Out & channel20_Kernel44_Valid_Out & channel21_Kernel44_Valid_Out & channel22_Kernel44_Valid_Out & channel23_Kernel44_Valid_Out & channel24_Kernel44_Valid_Out & channel25_Kernel44_Valid_Out & channel26_Kernel44_Valid_Out & channel27_Kernel44_Valid_Out & channel28_Kernel44_Valid_Out & channel29_Kernel44_Valid_Out & channel30_Kernel44_Valid_Out & channel31_Kernel44_Valid_Out & channel32_Kernel44_Valid_Out;

	wire channel1_Kernel45_Valid_Out, channel2_Kernel45_Valid_Out, channel3_Kernel45_Valid_Out, channel4_Kernel45_Valid_Out, channel5_Kernel45_Valid_Out, channel6_Kernel45_Valid_Out, channel7_Kernel45_Valid_Out, channel8_Kernel45_Valid_Out, channel9_Kernel45_Valid_Out, channel10_Kernel45_Valid_Out, channel11_Kernel45_Valid_Out, channel12_Kernel45_Valid_Out, channel13_Kernel45_Valid_Out, channel14_Kernel45_Valid_Out, channel15_Kernel45_Valid_Out, channel16_Kernel45_Valid_Out, channel17_Kernel45_Valid_Out, channel18_Kernel45_Valid_Out, channel19_Kernel45_Valid_Out, channel20_Kernel45_Valid_Out, channel21_Kernel45_Valid_Out, channel22_Kernel45_Valid_Out, channel23_Kernel45_Valid_Out, channel24_Kernel45_Valid_Out, channel25_Kernel45_Valid_Out, channel26_Kernel45_Valid_Out, channel27_Kernel45_Valid_Out, channel28_Kernel45_Valid_Out, channel29_Kernel45_Valid_Out, channel30_Kernel45_Valid_Out, channel31_Kernel45_Valid_Out, channel32_Kernel45_Valid_Out;

	assign add_kernel45=channel1_Kernel45_Valid_Out & channel2_Kernel45_Valid_Out & channel3_Kernel45_Valid_Out & channel4_Kernel45_Valid_Out & channel5_Kernel45_Valid_Out & channel6_Kernel45_Valid_Out & channel7_Kernel45_Valid_Out & channel8_Kernel45_Valid_Out & channel9_Kernel45_Valid_Out & channel10_Kernel45_Valid_Out & channel11_Kernel45_Valid_Out & channel12_Kernel45_Valid_Out & channel13_Kernel45_Valid_Out & channel14_Kernel45_Valid_Out & channel15_Kernel45_Valid_Out & channel16_Kernel45_Valid_Out & channel17_Kernel45_Valid_Out & channel18_Kernel45_Valid_Out & channel19_Kernel45_Valid_Out & channel20_Kernel45_Valid_Out & channel21_Kernel45_Valid_Out & channel22_Kernel45_Valid_Out & channel23_Kernel45_Valid_Out & channel24_Kernel45_Valid_Out & channel25_Kernel45_Valid_Out & channel26_Kernel45_Valid_Out & channel27_Kernel45_Valid_Out & channel28_Kernel45_Valid_Out & channel29_Kernel45_Valid_Out & channel30_Kernel45_Valid_Out & channel31_Kernel45_Valid_Out & channel32_Kernel45_Valid_Out;

	wire channel1_Kernel46_Valid_Out, channel2_Kernel46_Valid_Out, channel3_Kernel46_Valid_Out, channel4_Kernel46_Valid_Out, channel5_Kernel46_Valid_Out, channel6_Kernel46_Valid_Out, channel7_Kernel46_Valid_Out, channel8_Kernel46_Valid_Out, channel9_Kernel46_Valid_Out, channel10_Kernel46_Valid_Out, channel11_Kernel46_Valid_Out, channel12_Kernel46_Valid_Out, channel13_Kernel46_Valid_Out, channel14_Kernel46_Valid_Out, channel15_Kernel46_Valid_Out, channel16_Kernel46_Valid_Out, channel17_Kernel46_Valid_Out, channel18_Kernel46_Valid_Out, channel19_Kernel46_Valid_Out, channel20_Kernel46_Valid_Out, channel21_Kernel46_Valid_Out, channel22_Kernel46_Valid_Out, channel23_Kernel46_Valid_Out, channel24_Kernel46_Valid_Out, channel25_Kernel46_Valid_Out, channel26_Kernel46_Valid_Out, channel27_Kernel46_Valid_Out, channel28_Kernel46_Valid_Out, channel29_Kernel46_Valid_Out, channel30_Kernel46_Valid_Out, channel31_Kernel46_Valid_Out, channel32_Kernel46_Valid_Out;

	assign add_kernel46=channel1_Kernel46_Valid_Out & channel2_Kernel46_Valid_Out & channel3_Kernel46_Valid_Out & channel4_Kernel46_Valid_Out & channel5_Kernel46_Valid_Out & channel6_Kernel46_Valid_Out & channel7_Kernel46_Valid_Out & channel8_Kernel46_Valid_Out & channel9_Kernel46_Valid_Out & channel10_Kernel46_Valid_Out & channel11_Kernel46_Valid_Out & channel12_Kernel46_Valid_Out & channel13_Kernel46_Valid_Out & channel14_Kernel46_Valid_Out & channel15_Kernel46_Valid_Out & channel16_Kernel46_Valid_Out & channel17_Kernel46_Valid_Out & channel18_Kernel46_Valid_Out & channel19_Kernel46_Valid_Out & channel20_Kernel46_Valid_Out & channel21_Kernel46_Valid_Out & channel22_Kernel46_Valid_Out & channel23_Kernel46_Valid_Out & channel24_Kernel46_Valid_Out & channel25_Kernel46_Valid_Out & channel26_Kernel46_Valid_Out & channel27_Kernel46_Valid_Out & channel28_Kernel46_Valid_Out & channel29_Kernel46_Valid_Out & channel30_Kernel46_Valid_Out & channel31_Kernel46_Valid_Out & channel32_Kernel46_Valid_Out;

	wire channel1_Kernel47_Valid_Out, channel2_Kernel47_Valid_Out, channel3_Kernel47_Valid_Out, channel4_Kernel47_Valid_Out, channel5_Kernel47_Valid_Out, channel6_Kernel47_Valid_Out, channel7_Kernel47_Valid_Out, channel8_Kernel47_Valid_Out, channel9_Kernel47_Valid_Out, channel10_Kernel47_Valid_Out, channel11_Kernel47_Valid_Out, channel12_Kernel47_Valid_Out, channel13_Kernel47_Valid_Out, channel14_Kernel47_Valid_Out, channel15_Kernel47_Valid_Out, channel16_Kernel47_Valid_Out, channel17_Kernel47_Valid_Out, channel18_Kernel47_Valid_Out, channel19_Kernel47_Valid_Out, channel20_Kernel47_Valid_Out, channel21_Kernel47_Valid_Out, channel22_Kernel47_Valid_Out, channel23_Kernel47_Valid_Out, channel24_Kernel47_Valid_Out, channel25_Kernel47_Valid_Out, channel26_Kernel47_Valid_Out, channel27_Kernel47_Valid_Out, channel28_Kernel47_Valid_Out, channel29_Kernel47_Valid_Out, channel30_Kernel47_Valid_Out, channel31_Kernel47_Valid_Out, channel32_Kernel47_Valid_Out;

	assign add_kernel47=channel1_Kernel47_Valid_Out & channel2_Kernel47_Valid_Out & channel3_Kernel47_Valid_Out & channel4_Kernel47_Valid_Out & channel5_Kernel47_Valid_Out & channel6_Kernel47_Valid_Out & channel7_Kernel47_Valid_Out & channel8_Kernel47_Valid_Out & channel9_Kernel47_Valid_Out & channel10_Kernel47_Valid_Out & channel11_Kernel47_Valid_Out & channel12_Kernel47_Valid_Out & channel13_Kernel47_Valid_Out & channel14_Kernel47_Valid_Out & channel15_Kernel47_Valid_Out & channel16_Kernel47_Valid_Out & channel17_Kernel47_Valid_Out & channel18_Kernel47_Valid_Out & channel19_Kernel47_Valid_Out & channel20_Kernel47_Valid_Out & channel21_Kernel47_Valid_Out & channel22_Kernel47_Valid_Out & channel23_Kernel47_Valid_Out & channel24_Kernel47_Valid_Out & channel25_Kernel47_Valid_Out & channel26_Kernel47_Valid_Out & channel27_Kernel47_Valid_Out & channel28_Kernel47_Valid_Out & channel29_Kernel47_Valid_Out & channel30_Kernel47_Valid_Out & channel31_Kernel47_Valid_Out & channel32_Kernel47_Valid_Out;

	wire channel1_Kernel48_Valid_Out, channel2_Kernel48_Valid_Out, channel3_Kernel48_Valid_Out, channel4_Kernel48_Valid_Out, channel5_Kernel48_Valid_Out, channel6_Kernel48_Valid_Out, channel7_Kernel48_Valid_Out, channel8_Kernel48_Valid_Out, channel9_Kernel48_Valid_Out, channel10_Kernel48_Valid_Out, channel11_Kernel48_Valid_Out, channel12_Kernel48_Valid_Out, channel13_Kernel48_Valid_Out, channel14_Kernel48_Valid_Out, channel15_Kernel48_Valid_Out, channel16_Kernel48_Valid_Out, channel17_Kernel48_Valid_Out, channel18_Kernel48_Valid_Out, channel19_Kernel48_Valid_Out, channel20_Kernel48_Valid_Out, channel21_Kernel48_Valid_Out, channel22_Kernel48_Valid_Out, channel23_Kernel48_Valid_Out, channel24_Kernel48_Valid_Out, channel25_Kernel48_Valid_Out, channel26_Kernel48_Valid_Out, channel27_Kernel48_Valid_Out, channel28_Kernel48_Valid_Out, channel29_Kernel48_Valid_Out, channel30_Kernel48_Valid_Out, channel31_Kernel48_Valid_Out, channel32_Kernel48_Valid_Out;

	assign add_kernel48=channel1_Kernel48_Valid_Out & channel2_Kernel48_Valid_Out & channel3_Kernel48_Valid_Out & channel4_Kernel48_Valid_Out & channel5_Kernel48_Valid_Out & channel6_Kernel48_Valid_Out & channel7_Kernel48_Valid_Out & channel8_Kernel48_Valid_Out & channel9_Kernel48_Valid_Out & channel10_Kernel48_Valid_Out & channel11_Kernel48_Valid_Out & channel12_Kernel48_Valid_Out & channel13_Kernel48_Valid_Out & channel14_Kernel48_Valid_Out & channel15_Kernel48_Valid_Out & channel16_Kernel48_Valid_Out & channel17_Kernel48_Valid_Out & channel18_Kernel48_Valid_Out & channel19_Kernel48_Valid_Out & channel20_Kernel48_Valid_Out & channel21_Kernel48_Valid_Out & channel22_Kernel48_Valid_Out & channel23_Kernel48_Valid_Out & channel24_Kernel48_Valid_Out & channel25_Kernel48_Valid_Out & channel26_Kernel48_Valid_Out & channel27_Kernel48_Valid_Out & channel28_Kernel48_Valid_Out & channel29_Kernel48_Valid_Out & channel30_Kernel48_Valid_Out & channel31_Kernel48_Valid_Out & channel32_Kernel48_Valid_Out;

	wire channel1_Kernel49_Valid_Out, channel2_Kernel49_Valid_Out, channel3_Kernel49_Valid_Out, channel4_Kernel49_Valid_Out, channel5_Kernel49_Valid_Out, channel6_Kernel49_Valid_Out, channel7_Kernel49_Valid_Out, channel8_Kernel49_Valid_Out, channel9_Kernel49_Valid_Out, channel10_Kernel49_Valid_Out, channel11_Kernel49_Valid_Out, channel12_Kernel49_Valid_Out, channel13_Kernel49_Valid_Out, channel14_Kernel49_Valid_Out, channel15_Kernel49_Valid_Out, channel16_Kernel49_Valid_Out, channel17_Kernel49_Valid_Out, channel18_Kernel49_Valid_Out, channel19_Kernel49_Valid_Out, channel20_Kernel49_Valid_Out, channel21_Kernel49_Valid_Out, channel22_Kernel49_Valid_Out, channel23_Kernel49_Valid_Out, channel24_Kernel49_Valid_Out, channel25_Kernel49_Valid_Out, channel26_Kernel49_Valid_Out, channel27_Kernel49_Valid_Out, channel28_Kernel49_Valid_Out, channel29_Kernel49_Valid_Out, channel30_Kernel49_Valid_Out, channel31_Kernel49_Valid_Out, channel32_Kernel49_Valid_Out;

	assign add_kernel49=channel1_Kernel49_Valid_Out & channel2_Kernel49_Valid_Out & channel3_Kernel49_Valid_Out & channel4_Kernel49_Valid_Out & channel5_Kernel49_Valid_Out & channel6_Kernel49_Valid_Out & channel7_Kernel49_Valid_Out & channel8_Kernel49_Valid_Out & channel9_Kernel49_Valid_Out & channel10_Kernel49_Valid_Out & channel11_Kernel49_Valid_Out & channel12_Kernel49_Valid_Out & channel13_Kernel49_Valid_Out & channel14_Kernel49_Valid_Out & channel15_Kernel49_Valid_Out & channel16_Kernel49_Valid_Out & channel17_Kernel49_Valid_Out & channel18_Kernel49_Valid_Out & channel19_Kernel49_Valid_Out & channel20_Kernel49_Valid_Out & channel21_Kernel49_Valid_Out & channel22_Kernel49_Valid_Out & channel23_Kernel49_Valid_Out & channel24_Kernel49_Valid_Out & channel25_Kernel49_Valid_Out & channel26_Kernel49_Valid_Out & channel27_Kernel49_Valid_Out & channel28_Kernel49_Valid_Out & channel29_Kernel49_Valid_Out & channel30_Kernel49_Valid_Out & channel31_Kernel49_Valid_Out & channel32_Kernel49_Valid_Out;

	wire channel1_Kernel50_Valid_Out, channel2_Kernel50_Valid_Out, channel3_Kernel50_Valid_Out, channel4_Kernel50_Valid_Out, channel5_Kernel50_Valid_Out, channel6_Kernel50_Valid_Out, channel7_Kernel50_Valid_Out, channel8_Kernel50_Valid_Out, channel9_Kernel50_Valid_Out, channel10_Kernel50_Valid_Out, channel11_Kernel50_Valid_Out, channel12_Kernel50_Valid_Out, channel13_Kernel50_Valid_Out, channel14_Kernel50_Valid_Out, channel15_Kernel50_Valid_Out, channel16_Kernel50_Valid_Out, channel17_Kernel50_Valid_Out, channel18_Kernel50_Valid_Out, channel19_Kernel50_Valid_Out, channel20_Kernel50_Valid_Out, channel21_Kernel50_Valid_Out, channel22_Kernel50_Valid_Out, channel23_Kernel50_Valid_Out, channel24_Kernel50_Valid_Out, channel25_Kernel50_Valid_Out, channel26_Kernel50_Valid_Out, channel27_Kernel50_Valid_Out, channel28_Kernel50_Valid_Out, channel29_Kernel50_Valid_Out, channel30_Kernel50_Valid_Out, channel31_Kernel50_Valid_Out, channel32_Kernel50_Valid_Out;

	assign add_kernel50=channel1_Kernel50_Valid_Out & channel2_Kernel50_Valid_Out & channel3_Kernel50_Valid_Out & channel4_Kernel50_Valid_Out & channel5_Kernel50_Valid_Out & channel6_Kernel50_Valid_Out & channel7_Kernel50_Valid_Out & channel8_Kernel50_Valid_Out & channel9_Kernel50_Valid_Out & channel10_Kernel50_Valid_Out & channel11_Kernel50_Valid_Out & channel12_Kernel50_Valid_Out & channel13_Kernel50_Valid_Out & channel14_Kernel50_Valid_Out & channel15_Kernel50_Valid_Out & channel16_Kernel50_Valid_Out & channel17_Kernel50_Valid_Out & channel18_Kernel50_Valid_Out & channel19_Kernel50_Valid_Out & channel20_Kernel50_Valid_Out & channel21_Kernel50_Valid_Out & channel22_Kernel50_Valid_Out & channel23_Kernel50_Valid_Out & channel24_Kernel50_Valid_Out & channel25_Kernel50_Valid_Out & channel26_Kernel50_Valid_Out & channel27_Kernel50_Valid_Out & channel28_Kernel50_Valid_Out & channel29_Kernel50_Valid_Out & channel30_Kernel50_Valid_Out & channel31_Kernel50_Valid_Out & channel32_Kernel50_Valid_Out;

	wire channel1_Kernel51_Valid_Out, channel2_Kernel51_Valid_Out, channel3_Kernel51_Valid_Out, channel4_Kernel51_Valid_Out, channel5_Kernel51_Valid_Out, channel6_Kernel51_Valid_Out, channel7_Kernel51_Valid_Out, channel8_Kernel51_Valid_Out, channel9_Kernel51_Valid_Out, channel10_Kernel51_Valid_Out, channel11_Kernel51_Valid_Out, channel12_Kernel51_Valid_Out, channel13_Kernel51_Valid_Out, channel14_Kernel51_Valid_Out, channel15_Kernel51_Valid_Out, channel16_Kernel51_Valid_Out, channel17_Kernel51_Valid_Out, channel18_Kernel51_Valid_Out, channel19_Kernel51_Valid_Out, channel20_Kernel51_Valid_Out, channel21_Kernel51_Valid_Out, channel22_Kernel51_Valid_Out, channel23_Kernel51_Valid_Out, channel24_Kernel51_Valid_Out, channel25_Kernel51_Valid_Out, channel26_Kernel51_Valid_Out, channel27_Kernel51_Valid_Out, channel28_Kernel51_Valid_Out, channel29_Kernel51_Valid_Out, channel30_Kernel51_Valid_Out, channel31_Kernel51_Valid_Out, channel32_Kernel51_Valid_Out;

	assign add_kernel51=channel1_Kernel51_Valid_Out & channel2_Kernel51_Valid_Out & channel3_Kernel51_Valid_Out & channel4_Kernel51_Valid_Out & channel5_Kernel51_Valid_Out & channel6_Kernel51_Valid_Out & channel7_Kernel51_Valid_Out & channel8_Kernel51_Valid_Out & channel9_Kernel51_Valid_Out & channel10_Kernel51_Valid_Out & channel11_Kernel51_Valid_Out & channel12_Kernel51_Valid_Out & channel13_Kernel51_Valid_Out & channel14_Kernel51_Valid_Out & channel15_Kernel51_Valid_Out & channel16_Kernel51_Valid_Out & channel17_Kernel51_Valid_Out & channel18_Kernel51_Valid_Out & channel19_Kernel51_Valid_Out & channel20_Kernel51_Valid_Out & channel21_Kernel51_Valid_Out & channel22_Kernel51_Valid_Out & channel23_Kernel51_Valid_Out & channel24_Kernel51_Valid_Out & channel25_Kernel51_Valid_Out & channel26_Kernel51_Valid_Out & channel27_Kernel51_Valid_Out & channel28_Kernel51_Valid_Out & channel29_Kernel51_Valid_Out & channel30_Kernel51_Valid_Out & channel31_Kernel51_Valid_Out & channel32_Kernel51_Valid_Out;

	wire channel1_Kernel52_Valid_Out, channel2_Kernel52_Valid_Out, channel3_Kernel52_Valid_Out, channel4_Kernel52_Valid_Out, channel5_Kernel52_Valid_Out, channel6_Kernel52_Valid_Out, channel7_Kernel52_Valid_Out, channel8_Kernel52_Valid_Out, channel9_Kernel52_Valid_Out, channel10_Kernel52_Valid_Out, channel11_Kernel52_Valid_Out, channel12_Kernel52_Valid_Out, channel13_Kernel52_Valid_Out, channel14_Kernel52_Valid_Out, channel15_Kernel52_Valid_Out, channel16_Kernel52_Valid_Out, channel17_Kernel52_Valid_Out, channel18_Kernel52_Valid_Out, channel19_Kernel52_Valid_Out, channel20_Kernel52_Valid_Out, channel21_Kernel52_Valid_Out, channel22_Kernel52_Valid_Out, channel23_Kernel52_Valid_Out, channel24_Kernel52_Valid_Out, channel25_Kernel52_Valid_Out, channel26_Kernel52_Valid_Out, channel27_Kernel52_Valid_Out, channel28_Kernel52_Valid_Out, channel29_Kernel52_Valid_Out, channel30_Kernel52_Valid_Out, channel31_Kernel52_Valid_Out, channel32_Kernel52_Valid_Out;

	assign add_kernel52=channel1_Kernel52_Valid_Out & channel2_Kernel52_Valid_Out & channel3_Kernel52_Valid_Out & channel4_Kernel52_Valid_Out & channel5_Kernel52_Valid_Out & channel6_Kernel52_Valid_Out & channel7_Kernel52_Valid_Out & channel8_Kernel52_Valid_Out & channel9_Kernel52_Valid_Out & channel10_Kernel52_Valid_Out & channel11_Kernel52_Valid_Out & channel12_Kernel52_Valid_Out & channel13_Kernel52_Valid_Out & channel14_Kernel52_Valid_Out & channel15_Kernel52_Valid_Out & channel16_Kernel52_Valid_Out & channel17_Kernel52_Valid_Out & channel18_Kernel52_Valid_Out & channel19_Kernel52_Valid_Out & channel20_Kernel52_Valid_Out & channel21_Kernel52_Valid_Out & channel22_Kernel52_Valid_Out & channel23_Kernel52_Valid_Out & channel24_Kernel52_Valid_Out & channel25_Kernel52_Valid_Out & channel26_Kernel52_Valid_Out & channel27_Kernel52_Valid_Out & channel28_Kernel52_Valid_Out & channel29_Kernel52_Valid_Out & channel30_Kernel52_Valid_Out & channel31_Kernel52_Valid_Out & channel32_Kernel52_Valid_Out;

	wire channel1_Kernel53_Valid_Out, channel2_Kernel53_Valid_Out, channel3_Kernel53_Valid_Out, channel4_Kernel53_Valid_Out, channel5_Kernel53_Valid_Out, channel6_Kernel53_Valid_Out, channel7_Kernel53_Valid_Out, channel8_Kernel53_Valid_Out, channel9_Kernel53_Valid_Out, channel10_Kernel53_Valid_Out, channel11_Kernel53_Valid_Out, channel12_Kernel53_Valid_Out, channel13_Kernel53_Valid_Out, channel14_Kernel53_Valid_Out, channel15_Kernel53_Valid_Out, channel16_Kernel53_Valid_Out, channel17_Kernel53_Valid_Out, channel18_Kernel53_Valid_Out, channel19_Kernel53_Valid_Out, channel20_Kernel53_Valid_Out, channel21_Kernel53_Valid_Out, channel22_Kernel53_Valid_Out, channel23_Kernel53_Valid_Out, channel24_Kernel53_Valid_Out, channel25_Kernel53_Valid_Out, channel26_Kernel53_Valid_Out, channel27_Kernel53_Valid_Out, channel28_Kernel53_Valid_Out, channel29_Kernel53_Valid_Out, channel30_Kernel53_Valid_Out, channel31_Kernel53_Valid_Out, channel32_Kernel53_Valid_Out;

	assign add_kernel53=channel1_Kernel53_Valid_Out & channel2_Kernel53_Valid_Out & channel3_Kernel53_Valid_Out & channel4_Kernel53_Valid_Out & channel5_Kernel53_Valid_Out & channel6_Kernel53_Valid_Out & channel7_Kernel53_Valid_Out & channel8_Kernel53_Valid_Out & channel9_Kernel53_Valid_Out & channel10_Kernel53_Valid_Out & channel11_Kernel53_Valid_Out & channel12_Kernel53_Valid_Out & channel13_Kernel53_Valid_Out & channel14_Kernel53_Valid_Out & channel15_Kernel53_Valid_Out & channel16_Kernel53_Valid_Out & channel17_Kernel53_Valid_Out & channel18_Kernel53_Valid_Out & channel19_Kernel53_Valid_Out & channel20_Kernel53_Valid_Out & channel21_Kernel53_Valid_Out & channel22_Kernel53_Valid_Out & channel23_Kernel53_Valid_Out & channel24_Kernel53_Valid_Out & channel25_Kernel53_Valid_Out & channel26_Kernel53_Valid_Out & channel27_Kernel53_Valid_Out & channel28_Kernel53_Valid_Out & channel29_Kernel53_Valid_Out & channel30_Kernel53_Valid_Out & channel31_Kernel53_Valid_Out & channel32_Kernel53_Valid_Out;

	wire channel1_Kernel54_Valid_Out, channel2_Kernel54_Valid_Out, channel3_Kernel54_Valid_Out, channel4_Kernel54_Valid_Out, channel5_Kernel54_Valid_Out, channel6_Kernel54_Valid_Out, channel7_Kernel54_Valid_Out, channel8_Kernel54_Valid_Out, channel9_Kernel54_Valid_Out, channel10_Kernel54_Valid_Out, channel11_Kernel54_Valid_Out, channel12_Kernel54_Valid_Out, channel13_Kernel54_Valid_Out, channel14_Kernel54_Valid_Out, channel15_Kernel54_Valid_Out, channel16_Kernel54_Valid_Out, channel17_Kernel54_Valid_Out, channel18_Kernel54_Valid_Out, channel19_Kernel54_Valid_Out, channel20_Kernel54_Valid_Out, channel21_Kernel54_Valid_Out, channel22_Kernel54_Valid_Out, channel23_Kernel54_Valid_Out, channel24_Kernel54_Valid_Out, channel25_Kernel54_Valid_Out, channel26_Kernel54_Valid_Out, channel27_Kernel54_Valid_Out, channel28_Kernel54_Valid_Out, channel29_Kernel54_Valid_Out, channel30_Kernel54_Valid_Out, channel31_Kernel54_Valid_Out, channel32_Kernel54_Valid_Out;

	assign add_kernel54=channel1_Kernel54_Valid_Out & channel2_Kernel54_Valid_Out & channel3_Kernel54_Valid_Out & channel4_Kernel54_Valid_Out & channel5_Kernel54_Valid_Out & channel6_Kernel54_Valid_Out & channel7_Kernel54_Valid_Out & channel8_Kernel54_Valid_Out & channel9_Kernel54_Valid_Out & channel10_Kernel54_Valid_Out & channel11_Kernel54_Valid_Out & channel12_Kernel54_Valid_Out & channel13_Kernel54_Valid_Out & channel14_Kernel54_Valid_Out & channel15_Kernel54_Valid_Out & channel16_Kernel54_Valid_Out & channel17_Kernel54_Valid_Out & channel18_Kernel54_Valid_Out & channel19_Kernel54_Valid_Out & channel20_Kernel54_Valid_Out & channel21_Kernel54_Valid_Out & channel22_Kernel54_Valid_Out & channel23_Kernel54_Valid_Out & channel24_Kernel54_Valid_Out & channel25_Kernel54_Valid_Out & channel26_Kernel54_Valid_Out & channel27_Kernel54_Valid_Out & channel28_Kernel54_Valid_Out & channel29_Kernel54_Valid_Out & channel30_Kernel54_Valid_Out & channel31_Kernel54_Valid_Out & channel32_Kernel54_Valid_Out;

	wire channel1_Kernel55_Valid_Out, channel2_Kernel55_Valid_Out, channel3_Kernel55_Valid_Out, channel4_Kernel55_Valid_Out, channel5_Kernel55_Valid_Out, channel6_Kernel55_Valid_Out, channel7_Kernel55_Valid_Out, channel8_Kernel55_Valid_Out, channel9_Kernel55_Valid_Out, channel10_Kernel55_Valid_Out, channel11_Kernel55_Valid_Out, channel12_Kernel55_Valid_Out, channel13_Kernel55_Valid_Out, channel14_Kernel55_Valid_Out, channel15_Kernel55_Valid_Out, channel16_Kernel55_Valid_Out, channel17_Kernel55_Valid_Out, channel18_Kernel55_Valid_Out, channel19_Kernel55_Valid_Out, channel20_Kernel55_Valid_Out, channel21_Kernel55_Valid_Out, channel22_Kernel55_Valid_Out, channel23_Kernel55_Valid_Out, channel24_Kernel55_Valid_Out, channel25_Kernel55_Valid_Out, channel26_Kernel55_Valid_Out, channel27_Kernel55_Valid_Out, channel28_Kernel55_Valid_Out, channel29_Kernel55_Valid_Out, channel30_Kernel55_Valid_Out, channel31_Kernel55_Valid_Out, channel32_Kernel55_Valid_Out;

	assign add_kernel55=channel1_Kernel55_Valid_Out & channel2_Kernel55_Valid_Out & channel3_Kernel55_Valid_Out & channel4_Kernel55_Valid_Out & channel5_Kernel55_Valid_Out & channel6_Kernel55_Valid_Out & channel7_Kernel55_Valid_Out & channel8_Kernel55_Valid_Out & channel9_Kernel55_Valid_Out & channel10_Kernel55_Valid_Out & channel11_Kernel55_Valid_Out & channel12_Kernel55_Valid_Out & channel13_Kernel55_Valid_Out & channel14_Kernel55_Valid_Out & channel15_Kernel55_Valid_Out & channel16_Kernel55_Valid_Out & channel17_Kernel55_Valid_Out & channel18_Kernel55_Valid_Out & channel19_Kernel55_Valid_Out & channel20_Kernel55_Valid_Out & channel21_Kernel55_Valid_Out & channel22_Kernel55_Valid_Out & channel23_Kernel55_Valid_Out & channel24_Kernel55_Valid_Out & channel25_Kernel55_Valid_Out & channel26_Kernel55_Valid_Out & channel27_Kernel55_Valid_Out & channel28_Kernel55_Valid_Out & channel29_Kernel55_Valid_Out & channel30_Kernel55_Valid_Out & channel31_Kernel55_Valid_Out & channel32_Kernel55_Valid_Out;

	wire channel1_Kernel56_Valid_Out, channel2_Kernel56_Valid_Out, channel3_Kernel56_Valid_Out, channel4_Kernel56_Valid_Out, channel5_Kernel56_Valid_Out, channel6_Kernel56_Valid_Out, channel7_Kernel56_Valid_Out, channel8_Kernel56_Valid_Out, channel9_Kernel56_Valid_Out, channel10_Kernel56_Valid_Out, channel11_Kernel56_Valid_Out, channel12_Kernel56_Valid_Out, channel13_Kernel56_Valid_Out, channel14_Kernel56_Valid_Out, channel15_Kernel56_Valid_Out, channel16_Kernel56_Valid_Out, channel17_Kernel56_Valid_Out, channel18_Kernel56_Valid_Out, channel19_Kernel56_Valid_Out, channel20_Kernel56_Valid_Out, channel21_Kernel56_Valid_Out, channel22_Kernel56_Valid_Out, channel23_Kernel56_Valid_Out, channel24_Kernel56_Valid_Out, channel25_Kernel56_Valid_Out, channel26_Kernel56_Valid_Out, channel27_Kernel56_Valid_Out, channel28_Kernel56_Valid_Out, channel29_Kernel56_Valid_Out, channel30_Kernel56_Valid_Out, channel31_Kernel56_Valid_Out, channel32_Kernel56_Valid_Out;

	assign add_kernel56=channel1_Kernel56_Valid_Out & channel2_Kernel56_Valid_Out & channel3_Kernel56_Valid_Out & channel4_Kernel56_Valid_Out & channel5_Kernel56_Valid_Out & channel6_Kernel56_Valid_Out & channel7_Kernel56_Valid_Out & channel8_Kernel56_Valid_Out & channel9_Kernel56_Valid_Out & channel10_Kernel56_Valid_Out & channel11_Kernel56_Valid_Out & channel12_Kernel56_Valid_Out & channel13_Kernel56_Valid_Out & channel14_Kernel56_Valid_Out & channel15_Kernel56_Valid_Out & channel16_Kernel56_Valid_Out & channel17_Kernel56_Valid_Out & channel18_Kernel56_Valid_Out & channel19_Kernel56_Valid_Out & channel20_Kernel56_Valid_Out & channel21_Kernel56_Valid_Out & channel22_Kernel56_Valid_Out & channel23_Kernel56_Valid_Out & channel24_Kernel56_Valid_Out & channel25_Kernel56_Valid_Out & channel26_Kernel56_Valid_Out & channel27_Kernel56_Valid_Out & channel28_Kernel56_Valid_Out & channel29_Kernel56_Valid_Out & channel30_Kernel56_Valid_Out & channel31_Kernel56_Valid_Out & channel32_Kernel56_Valid_Out;

	wire channel1_Kernel57_Valid_Out, channel2_Kernel57_Valid_Out, channel3_Kernel57_Valid_Out, channel4_Kernel57_Valid_Out, channel5_Kernel57_Valid_Out, channel6_Kernel57_Valid_Out, channel7_Kernel57_Valid_Out, channel8_Kernel57_Valid_Out, channel9_Kernel57_Valid_Out, channel10_Kernel57_Valid_Out, channel11_Kernel57_Valid_Out, channel12_Kernel57_Valid_Out, channel13_Kernel57_Valid_Out, channel14_Kernel57_Valid_Out, channel15_Kernel57_Valid_Out, channel16_Kernel57_Valid_Out, channel17_Kernel57_Valid_Out, channel18_Kernel57_Valid_Out, channel19_Kernel57_Valid_Out, channel20_Kernel57_Valid_Out, channel21_Kernel57_Valid_Out, channel22_Kernel57_Valid_Out, channel23_Kernel57_Valid_Out, channel24_Kernel57_Valid_Out, channel25_Kernel57_Valid_Out, channel26_Kernel57_Valid_Out, channel27_Kernel57_Valid_Out, channel28_Kernel57_Valid_Out, channel29_Kernel57_Valid_Out, channel30_Kernel57_Valid_Out, channel31_Kernel57_Valid_Out, channel32_Kernel57_Valid_Out;

	assign add_kernel57=channel1_Kernel57_Valid_Out & channel2_Kernel57_Valid_Out & channel3_Kernel57_Valid_Out & channel4_Kernel57_Valid_Out & channel5_Kernel57_Valid_Out & channel6_Kernel57_Valid_Out & channel7_Kernel57_Valid_Out & channel8_Kernel57_Valid_Out & channel9_Kernel57_Valid_Out & channel10_Kernel57_Valid_Out & channel11_Kernel57_Valid_Out & channel12_Kernel57_Valid_Out & channel13_Kernel57_Valid_Out & channel14_Kernel57_Valid_Out & channel15_Kernel57_Valid_Out & channel16_Kernel57_Valid_Out & channel17_Kernel57_Valid_Out & channel18_Kernel57_Valid_Out & channel19_Kernel57_Valid_Out & channel20_Kernel57_Valid_Out & channel21_Kernel57_Valid_Out & channel22_Kernel57_Valid_Out & channel23_Kernel57_Valid_Out & channel24_Kernel57_Valid_Out & channel25_Kernel57_Valid_Out & channel26_Kernel57_Valid_Out & channel27_Kernel57_Valid_Out & channel28_Kernel57_Valid_Out & channel29_Kernel57_Valid_Out & channel30_Kernel57_Valid_Out & channel31_Kernel57_Valid_Out & channel32_Kernel57_Valid_Out;

	wire channel1_Kernel58_Valid_Out, channel2_Kernel58_Valid_Out, channel3_Kernel58_Valid_Out, channel4_Kernel58_Valid_Out, channel5_Kernel58_Valid_Out, channel6_Kernel58_Valid_Out, channel7_Kernel58_Valid_Out, channel8_Kernel58_Valid_Out, channel9_Kernel58_Valid_Out, channel10_Kernel58_Valid_Out, channel11_Kernel58_Valid_Out, channel12_Kernel58_Valid_Out, channel13_Kernel58_Valid_Out, channel14_Kernel58_Valid_Out, channel15_Kernel58_Valid_Out, channel16_Kernel58_Valid_Out, channel17_Kernel58_Valid_Out, channel18_Kernel58_Valid_Out, channel19_Kernel58_Valid_Out, channel20_Kernel58_Valid_Out, channel21_Kernel58_Valid_Out, channel22_Kernel58_Valid_Out, channel23_Kernel58_Valid_Out, channel24_Kernel58_Valid_Out, channel25_Kernel58_Valid_Out, channel26_Kernel58_Valid_Out, channel27_Kernel58_Valid_Out, channel28_Kernel58_Valid_Out, channel29_Kernel58_Valid_Out, channel30_Kernel58_Valid_Out, channel31_Kernel58_Valid_Out, channel32_Kernel58_Valid_Out;

	assign add_kernel58=channel1_Kernel58_Valid_Out & channel2_Kernel58_Valid_Out & channel3_Kernel58_Valid_Out & channel4_Kernel58_Valid_Out & channel5_Kernel58_Valid_Out & channel6_Kernel58_Valid_Out & channel7_Kernel58_Valid_Out & channel8_Kernel58_Valid_Out & channel9_Kernel58_Valid_Out & channel10_Kernel58_Valid_Out & channel11_Kernel58_Valid_Out & channel12_Kernel58_Valid_Out & channel13_Kernel58_Valid_Out & channel14_Kernel58_Valid_Out & channel15_Kernel58_Valid_Out & channel16_Kernel58_Valid_Out & channel17_Kernel58_Valid_Out & channel18_Kernel58_Valid_Out & channel19_Kernel58_Valid_Out & channel20_Kernel58_Valid_Out & channel21_Kernel58_Valid_Out & channel22_Kernel58_Valid_Out & channel23_Kernel58_Valid_Out & channel24_Kernel58_Valid_Out & channel25_Kernel58_Valid_Out & channel26_Kernel58_Valid_Out & channel27_Kernel58_Valid_Out & channel28_Kernel58_Valid_Out & channel29_Kernel58_Valid_Out & channel30_Kernel58_Valid_Out & channel31_Kernel58_Valid_Out & channel32_Kernel58_Valid_Out;

	wire channel1_Kernel59_Valid_Out, channel2_Kernel59_Valid_Out, channel3_Kernel59_Valid_Out, channel4_Kernel59_Valid_Out, channel5_Kernel59_Valid_Out, channel6_Kernel59_Valid_Out, channel7_Kernel59_Valid_Out, channel8_Kernel59_Valid_Out, channel9_Kernel59_Valid_Out, channel10_Kernel59_Valid_Out, channel11_Kernel59_Valid_Out, channel12_Kernel59_Valid_Out, channel13_Kernel59_Valid_Out, channel14_Kernel59_Valid_Out, channel15_Kernel59_Valid_Out, channel16_Kernel59_Valid_Out, channel17_Kernel59_Valid_Out, channel18_Kernel59_Valid_Out, channel19_Kernel59_Valid_Out, channel20_Kernel59_Valid_Out, channel21_Kernel59_Valid_Out, channel22_Kernel59_Valid_Out, channel23_Kernel59_Valid_Out, channel24_Kernel59_Valid_Out, channel25_Kernel59_Valid_Out, channel26_Kernel59_Valid_Out, channel27_Kernel59_Valid_Out, channel28_Kernel59_Valid_Out, channel29_Kernel59_Valid_Out, channel30_Kernel59_Valid_Out, channel31_Kernel59_Valid_Out, channel32_Kernel59_Valid_Out;

	assign add_kernel59=channel1_Kernel59_Valid_Out & channel2_Kernel59_Valid_Out & channel3_Kernel59_Valid_Out & channel4_Kernel59_Valid_Out & channel5_Kernel59_Valid_Out & channel6_Kernel59_Valid_Out & channel7_Kernel59_Valid_Out & channel8_Kernel59_Valid_Out & channel9_Kernel59_Valid_Out & channel10_Kernel59_Valid_Out & channel11_Kernel59_Valid_Out & channel12_Kernel59_Valid_Out & channel13_Kernel59_Valid_Out & channel14_Kernel59_Valid_Out & channel15_Kernel59_Valid_Out & channel16_Kernel59_Valid_Out & channel17_Kernel59_Valid_Out & channel18_Kernel59_Valid_Out & channel19_Kernel59_Valid_Out & channel20_Kernel59_Valid_Out & channel21_Kernel59_Valid_Out & channel22_Kernel59_Valid_Out & channel23_Kernel59_Valid_Out & channel24_Kernel59_Valid_Out & channel25_Kernel59_Valid_Out & channel26_Kernel59_Valid_Out & channel27_Kernel59_Valid_Out & channel28_Kernel59_Valid_Out & channel29_Kernel59_Valid_Out & channel30_Kernel59_Valid_Out & channel31_Kernel59_Valid_Out & channel32_Kernel59_Valid_Out;

	wire channel1_Kernel60_Valid_Out, channel2_Kernel60_Valid_Out, channel3_Kernel60_Valid_Out, channel4_Kernel60_Valid_Out, channel5_Kernel60_Valid_Out, channel6_Kernel60_Valid_Out, channel7_Kernel60_Valid_Out, channel8_Kernel60_Valid_Out, channel9_Kernel60_Valid_Out, channel10_Kernel60_Valid_Out, channel11_Kernel60_Valid_Out, channel12_Kernel60_Valid_Out, channel13_Kernel60_Valid_Out, channel14_Kernel60_Valid_Out, channel15_Kernel60_Valid_Out, channel16_Kernel60_Valid_Out, channel17_Kernel60_Valid_Out, channel18_Kernel60_Valid_Out, channel19_Kernel60_Valid_Out, channel20_Kernel60_Valid_Out, channel21_Kernel60_Valid_Out, channel22_Kernel60_Valid_Out, channel23_Kernel60_Valid_Out, channel24_Kernel60_Valid_Out, channel25_Kernel60_Valid_Out, channel26_Kernel60_Valid_Out, channel27_Kernel60_Valid_Out, channel28_Kernel60_Valid_Out, channel29_Kernel60_Valid_Out, channel30_Kernel60_Valid_Out, channel31_Kernel60_Valid_Out, channel32_Kernel60_Valid_Out;

	assign add_kernel60=channel1_Kernel60_Valid_Out & channel2_Kernel60_Valid_Out & channel3_Kernel60_Valid_Out & channel4_Kernel60_Valid_Out & channel5_Kernel60_Valid_Out & channel6_Kernel60_Valid_Out & channel7_Kernel60_Valid_Out & channel8_Kernel60_Valid_Out & channel9_Kernel60_Valid_Out & channel10_Kernel60_Valid_Out & channel11_Kernel60_Valid_Out & channel12_Kernel60_Valid_Out & channel13_Kernel60_Valid_Out & channel14_Kernel60_Valid_Out & channel15_Kernel60_Valid_Out & channel16_Kernel60_Valid_Out & channel17_Kernel60_Valid_Out & channel18_Kernel60_Valid_Out & channel19_Kernel60_Valid_Out & channel20_Kernel60_Valid_Out & channel21_Kernel60_Valid_Out & channel22_Kernel60_Valid_Out & channel23_Kernel60_Valid_Out & channel24_Kernel60_Valid_Out & channel25_Kernel60_Valid_Out & channel26_Kernel60_Valid_Out & channel27_Kernel60_Valid_Out & channel28_Kernel60_Valid_Out & channel29_Kernel60_Valid_Out & channel30_Kernel60_Valid_Out & channel31_Kernel60_Valid_Out & channel32_Kernel60_Valid_Out;

	wire channel1_Kernel61_Valid_Out, channel2_Kernel61_Valid_Out, channel3_Kernel61_Valid_Out, channel4_Kernel61_Valid_Out, channel5_Kernel61_Valid_Out, channel6_Kernel61_Valid_Out, channel7_Kernel61_Valid_Out, channel8_Kernel61_Valid_Out, channel9_Kernel61_Valid_Out, channel10_Kernel61_Valid_Out, channel11_Kernel61_Valid_Out, channel12_Kernel61_Valid_Out, channel13_Kernel61_Valid_Out, channel14_Kernel61_Valid_Out, channel15_Kernel61_Valid_Out, channel16_Kernel61_Valid_Out, channel17_Kernel61_Valid_Out, channel18_Kernel61_Valid_Out, channel19_Kernel61_Valid_Out, channel20_Kernel61_Valid_Out, channel21_Kernel61_Valid_Out, channel22_Kernel61_Valid_Out, channel23_Kernel61_Valid_Out, channel24_Kernel61_Valid_Out, channel25_Kernel61_Valid_Out, channel26_Kernel61_Valid_Out, channel27_Kernel61_Valid_Out, channel28_Kernel61_Valid_Out, channel29_Kernel61_Valid_Out, channel30_Kernel61_Valid_Out, channel31_Kernel61_Valid_Out, channel32_Kernel61_Valid_Out;

	assign add_kernel61=channel1_Kernel61_Valid_Out & channel2_Kernel61_Valid_Out & channel3_Kernel61_Valid_Out & channel4_Kernel61_Valid_Out & channel5_Kernel61_Valid_Out & channel6_Kernel61_Valid_Out & channel7_Kernel61_Valid_Out & channel8_Kernel61_Valid_Out & channel9_Kernel61_Valid_Out & channel10_Kernel61_Valid_Out & channel11_Kernel61_Valid_Out & channel12_Kernel61_Valid_Out & channel13_Kernel61_Valid_Out & channel14_Kernel61_Valid_Out & channel15_Kernel61_Valid_Out & channel16_Kernel61_Valid_Out & channel17_Kernel61_Valid_Out & channel18_Kernel61_Valid_Out & channel19_Kernel61_Valid_Out & channel20_Kernel61_Valid_Out & channel21_Kernel61_Valid_Out & channel22_Kernel61_Valid_Out & channel23_Kernel61_Valid_Out & channel24_Kernel61_Valid_Out & channel25_Kernel61_Valid_Out & channel26_Kernel61_Valid_Out & channel27_Kernel61_Valid_Out & channel28_Kernel61_Valid_Out & channel29_Kernel61_Valid_Out & channel30_Kernel61_Valid_Out & channel31_Kernel61_Valid_Out & channel32_Kernel61_Valid_Out;

	wire channel1_Kernel62_Valid_Out, channel2_Kernel62_Valid_Out, channel3_Kernel62_Valid_Out, channel4_Kernel62_Valid_Out, channel5_Kernel62_Valid_Out, channel6_Kernel62_Valid_Out, channel7_Kernel62_Valid_Out, channel8_Kernel62_Valid_Out, channel9_Kernel62_Valid_Out, channel10_Kernel62_Valid_Out, channel11_Kernel62_Valid_Out, channel12_Kernel62_Valid_Out, channel13_Kernel62_Valid_Out, channel14_Kernel62_Valid_Out, channel15_Kernel62_Valid_Out, channel16_Kernel62_Valid_Out, channel17_Kernel62_Valid_Out, channel18_Kernel62_Valid_Out, channel19_Kernel62_Valid_Out, channel20_Kernel62_Valid_Out, channel21_Kernel62_Valid_Out, channel22_Kernel62_Valid_Out, channel23_Kernel62_Valid_Out, channel24_Kernel62_Valid_Out, channel25_Kernel62_Valid_Out, channel26_Kernel62_Valid_Out, channel27_Kernel62_Valid_Out, channel28_Kernel62_Valid_Out, channel29_Kernel62_Valid_Out, channel30_Kernel62_Valid_Out, channel31_Kernel62_Valid_Out, channel32_Kernel62_Valid_Out;

	assign add_kernel62=channel1_Kernel62_Valid_Out & channel2_Kernel62_Valid_Out & channel3_Kernel62_Valid_Out & channel4_Kernel62_Valid_Out & channel5_Kernel62_Valid_Out & channel6_Kernel62_Valid_Out & channel7_Kernel62_Valid_Out & channel8_Kernel62_Valid_Out & channel9_Kernel62_Valid_Out & channel10_Kernel62_Valid_Out & channel11_Kernel62_Valid_Out & channel12_Kernel62_Valid_Out & channel13_Kernel62_Valid_Out & channel14_Kernel62_Valid_Out & channel15_Kernel62_Valid_Out & channel16_Kernel62_Valid_Out & channel17_Kernel62_Valid_Out & channel18_Kernel62_Valid_Out & channel19_Kernel62_Valid_Out & channel20_Kernel62_Valid_Out & channel21_Kernel62_Valid_Out & channel22_Kernel62_Valid_Out & channel23_Kernel62_Valid_Out & channel24_Kernel62_Valid_Out & channel25_Kernel62_Valid_Out & channel26_Kernel62_Valid_Out & channel27_Kernel62_Valid_Out & channel28_Kernel62_Valid_Out & channel29_Kernel62_Valid_Out & channel30_Kernel62_Valid_Out & channel31_Kernel62_Valid_Out & channel32_Kernel62_Valid_Out;

	wire channel1_Kernel63_Valid_Out, channel2_Kernel63_Valid_Out, channel3_Kernel63_Valid_Out, channel4_Kernel63_Valid_Out, channel5_Kernel63_Valid_Out, channel6_Kernel63_Valid_Out, channel7_Kernel63_Valid_Out, channel8_Kernel63_Valid_Out, channel9_Kernel63_Valid_Out, channel10_Kernel63_Valid_Out, channel11_Kernel63_Valid_Out, channel12_Kernel63_Valid_Out, channel13_Kernel63_Valid_Out, channel14_Kernel63_Valid_Out, channel15_Kernel63_Valid_Out, channel16_Kernel63_Valid_Out, channel17_Kernel63_Valid_Out, channel18_Kernel63_Valid_Out, channel19_Kernel63_Valid_Out, channel20_Kernel63_Valid_Out, channel21_Kernel63_Valid_Out, channel22_Kernel63_Valid_Out, channel23_Kernel63_Valid_Out, channel24_Kernel63_Valid_Out, channel25_Kernel63_Valid_Out, channel26_Kernel63_Valid_Out, channel27_Kernel63_Valid_Out, channel28_Kernel63_Valid_Out, channel29_Kernel63_Valid_Out, channel30_Kernel63_Valid_Out, channel31_Kernel63_Valid_Out, channel32_Kernel63_Valid_Out;

	assign add_kernel63=channel1_Kernel63_Valid_Out & channel2_Kernel63_Valid_Out & channel3_Kernel63_Valid_Out & channel4_Kernel63_Valid_Out & channel5_Kernel63_Valid_Out & channel6_Kernel63_Valid_Out & channel7_Kernel63_Valid_Out & channel8_Kernel63_Valid_Out & channel9_Kernel63_Valid_Out & channel10_Kernel63_Valid_Out & channel11_Kernel63_Valid_Out & channel12_Kernel63_Valid_Out & channel13_Kernel63_Valid_Out & channel14_Kernel63_Valid_Out & channel15_Kernel63_Valid_Out & channel16_Kernel63_Valid_Out & channel17_Kernel63_Valid_Out & channel18_Kernel63_Valid_Out & channel19_Kernel63_Valid_Out & channel20_Kernel63_Valid_Out & channel21_Kernel63_Valid_Out & channel22_Kernel63_Valid_Out & channel23_Kernel63_Valid_Out & channel24_Kernel63_Valid_Out & channel25_Kernel63_Valid_Out & channel26_Kernel63_Valid_Out & channel27_Kernel63_Valid_Out & channel28_Kernel63_Valid_Out & channel29_Kernel63_Valid_Out & channel30_Kernel63_Valid_Out & channel31_Kernel63_Valid_Out & channel32_Kernel63_Valid_Out;

	wire channel1_Kernel64_Valid_Out, channel2_Kernel64_Valid_Out, channel3_Kernel64_Valid_Out, channel4_Kernel64_Valid_Out, channel5_Kernel64_Valid_Out, channel6_Kernel64_Valid_Out, channel7_Kernel64_Valid_Out, channel8_Kernel64_Valid_Out, channel9_Kernel64_Valid_Out, channel10_Kernel64_Valid_Out, channel11_Kernel64_Valid_Out, channel12_Kernel64_Valid_Out, channel13_Kernel64_Valid_Out, channel14_Kernel64_Valid_Out, channel15_Kernel64_Valid_Out, channel16_Kernel64_Valid_Out, channel17_Kernel64_Valid_Out, channel18_Kernel64_Valid_Out, channel19_Kernel64_Valid_Out, channel20_Kernel64_Valid_Out, channel21_Kernel64_Valid_Out, channel22_Kernel64_Valid_Out, channel23_Kernel64_Valid_Out, channel24_Kernel64_Valid_Out, channel25_Kernel64_Valid_Out, channel26_Kernel64_Valid_Out, channel27_Kernel64_Valid_Out, channel28_Kernel64_Valid_Out, channel29_Kernel64_Valid_Out, channel30_Kernel64_Valid_Out, channel31_Kernel64_Valid_Out, channel32_Kernel64_Valid_Out;

	assign add_kernel64=channel1_Kernel64_Valid_Out & channel2_Kernel64_Valid_Out & channel3_Kernel64_Valid_Out & channel4_Kernel64_Valid_Out & channel5_Kernel64_Valid_Out & channel6_Kernel64_Valid_Out & channel7_Kernel64_Valid_Out & channel8_Kernel64_Valid_Out & channel9_Kernel64_Valid_Out & channel10_Kernel64_Valid_Out & channel11_Kernel64_Valid_Out & channel12_Kernel64_Valid_Out & channel13_Kernel64_Valid_Out & channel14_Kernel64_Valid_Out & channel15_Kernel64_Valid_Out & channel16_Kernel64_Valid_Out & channel17_Kernel64_Valid_Out & channel18_Kernel64_Valid_Out & channel19_Kernel64_Valid_Out & channel20_Kernel64_Valid_Out & channel21_Kernel64_Valid_Out & channel22_Kernel64_Valid_Out & channel23_Kernel64_Valid_Out & channel24_Kernel64_Valid_Out & channel25_Kernel64_Valid_Out & channel26_Kernel64_Valid_Out & channel27_Kernel64_Valid_Out & channel28_Kernel64_Valid_Out & channel29_Kernel64_Valid_Out & channel30_Kernel64_Valid_Out & channel31_Kernel64_Valid_Out & channel32_Kernel64_Valid_Out;


	wire [31:0] bn1_Data_Out, bn2_Data_Out, bn3_Data_Out, bn4_Data_Out, bn5_Data_Out, bn6_Data_Out, bn7_Data_Out, bn8_Data_Out, bn9_Data_Out, bn10_Data_Out, bn11_Data_Out, bn12_Data_Out, bn13_Data_Out, bn14_Data_Out, bn15_Data_Out, bn16_Data_Out, bn17_Data_Out, bn18_Data_Out, bn19_Data_Out, bn20_Data_Out, bn21_Data_Out, bn22_Data_Out, bn23_Data_Out, bn24_Data_Out, bn25_Data_Out, bn26_Data_Out, bn27_Data_Out, bn28_Data_Out, bn29_Data_Out, bn30_Data_Out, bn31_Data_Out, bn32_Data_Out, bn33_Data_Out, bn34_Data_Out, bn35_Data_Out, bn36_Data_Out, bn37_Data_Out, bn38_Data_Out, bn39_Data_Out, bn40_Data_Out, bn41_Data_Out, bn42_Data_Out, bn43_Data_Out, bn44_Data_Out, bn45_Data_Out, bn46_Data_Out, bn47_Data_Out, bn48_Data_Out, bn49_Data_Out, bn50_Data_Out, bn51_Data_Out, bn52_Data_Out, bn53_Data_Out, bn54_Data_Out, bn55_Data_Out, bn56_Data_Out, bn57_Data_Out, bn58_Data_Out, bn59_Data_Out, bn60_Data_Out, bn61_Data_Out, bn62_Data_Out, bn63_Data_Out, bn64_Data_Out;

	wire bn1_Valid_Out, bn2_Valid_Out, bn3_Valid_Out, bn4_Valid_Out, bn5_Valid_Out, bn6_Valid_Out, bn7_Valid_Out, bn8_Valid_Out, bn9_Valid_Out, bn10_Valid_Out, bn11_Valid_Out, bn12_Valid_Out, bn13_Valid_Out, bn14_Valid_Out, bn15_Valid_Out, bn16_Valid_Out, bn17_Valid_Out, bn18_Valid_Out, bn19_Valid_Out, bn20_Valid_Out, bn21_Valid_Out, bn22_Valid_Out, bn23_Valid_Out, bn24_Valid_Out, bn25_Valid_Out, bn26_Valid_Out, bn27_Valid_Out, bn28_Valid_Out, bn29_Valid_Out, bn30_Valid_Out, bn31_Valid_Out, bn32_Valid_Out, bn33_Valid_Out, bn34_Valid_Out, bn35_Valid_Out, bn36_Valid_Out, bn37_Valid_Out, bn38_Valid_Out, bn39_Valid_Out, bn40_Valid_Out, bn41_Valid_Out, bn42_Valid_Out, bn43_Valid_Out, bn44_Valid_Out, bn45_Valid_Out, bn46_Valid_Out, bn47_Valid_Out, bn48_Valid_Out, bn49_Valid_Out, bn50_Valid_Out, bn51_Valid_Out, bn52_Valid_Out, bn53_Valid_Out, bn54_Valid_Out, bn55_Valid_Out, bn56_Valid_Out, bn57_Valid_Out, bn58_Valid_Out, bn59_Valid_Out, bn60_Valid_Out, bn61_Valid_Out, bn62_Valid_Out, bn63_Valid_Out, bn64_Valid_Out;

	wire rl1_Valid_Out, rl2_Valid_Out, rl3_Valid_Out, rl4_Valid_Out, rl5_Valid_Out, rl6_Valid_Out, rl7_Valid_Out, rl8_Valid_Out, rl9_Valid_Out, rl10_Valid_Out, rl11_Valid_Out, rl12_Valid_Out, rl13_Valid_Out, rl14_Valid_Out, rl15_Valid_Out, rl16_Valid_Out, rl17_Valid_Out, rl18_Valid_Out, rl19_Valid_Out, rl20_Valid_Out, rl21_Valid_Out, rl22_Valid_Out, rl23_Valid_Out, rl24_Valid_Out, rl25_Valid_Out, rl26_Valid_Out, rl27_Valid_Out, rl28_Valid_Out, rl29_Valid_Out, rl30_Valid_Out, rl31_Valid_Out, rl32_Valid_Out, rl33_Valid_Out, rl34_Valid_Out, rl35_Valid_Out, rl36_Valid_Out, rl37_Valid_Out, rl38_Valid_Out, rl39_Valid_Out, rl40_Valid_Out, rl41_Valid_Out, rl42_Valid_Out, rl43_Valid_Out, rl44_Valid_Out, rl45_Valid_Out, rl46_Valid_Out, rl47_Valid_Out, rl48_Valid_Out, rl49_Valid_Out, rl50_Valid_Out, rl51_Valid_Out, rl52_Valid_Out, rl53_Valid_Out, rl54_Valid_Out, rl55_Valid_Out, rl56_Valid_Out, rl57_Valid_Out, rl58_Valid_Out, rl59_Valid_Out, rl60_Valid_Out, rl61_Valid_Out, rl62_Valid_Out, rl63_Valid_Out, rl64_Valid_Out;

	 assign Valid_Out = rl1_Valid_Out & rl2_Valid_Out & rl3_Valid_Out & rl4_Valid_Out & rl5_Valid_Out & rl6_Valid_Out & rl7_Valid_Out & rl8_Valid_Out & rl9_Valid_Out & rl10_Valid_Out & rl11_Valid_Out & rl12_Valid_Out & rl13_Valid_Out & rl14_Valid_Out & rl15_Valid_Out & rl16_Valid_Out & rl17_Valid_Out & rl18_Valid_Out & rl19_Valid_Out & rl20_Valid_Out & rl21_Valid_Out & rl22_Valid_Out & rl23_Valid_Out & rl24_Valid_Out & rl25_Valid_Out & rl26_Valid_Out & rl27_Valid_Out & rl28_Valid_Out & rl29_Valid_Out & rl30_Valid_Out & rl31_Valid_Out & rl32_Valid_Out & rl33_Valid_Out & rl34_Valid_Out & rl35_Valid_Out & rl36_Valid_Out & rl37_Valid_Out & rl38_Valid_Out & rl39_Valid_Out & rl40_Valid_Out & rl41_Valid_Out & rl42_Valid_Out & rl43_Valid_Out & rl44_Valid_Out & rl45_Valid_Out & rl46_Valid_Out & rl47_Valid_Out & rl48_Valid_Out & rl49_Valid_Out & rl50_Valid_Out & rl51_Valid_Out & rl52_Valid_Out & rl53_Valid_Out & rl54_Valid_Out & rl55_Valid_Out & rl56_Valid_Out & rl57_Valid_Out & rl58_Valid_Out & rl59_Valid_Out & rl60_Valid_Out & rl61_Valid_Out & rl62_Valid_Out & rl63_Valid_Out & rl64_Valid_Out;
//////////KERNEL1//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111101101110010001100010000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110011101100000101000000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110010011010111101101000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110001101000100110100110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111110100011001000110001010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111101110100000100111101101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111101110111100010110011011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111110111001111011101110110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110110010011010100111001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111101100010011100100110100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111111000011000011000001101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110010100001010010000110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111101001100001110111110100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111110011101011111000000001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111101110101001011110000000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111110011101001001100010110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111110011001000000000101100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111111010000111010000100001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111111011000000111101000011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111111000011011101110000000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111101011011100010100111001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111111010110000011101111001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111111000001111110001100011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111101001110101101001000111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111110110001111011100010000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110010100111010111110010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111101000001001100101010010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111110001001010001110011110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111110000101111011001100101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111111000111000000001111111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111110001010011110111000011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111101100011011101010010100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel1_Valid_Out)
	);
	Adder_32input add_k1(
		.Data1(Data_Out_Kernel1[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel1[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel1[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel1[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel1[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel1[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel1[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel1[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel1[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel1[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel1[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel1[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel1[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel1[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel1[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel1[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel1[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel1[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel1[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel1[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel1[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel1[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel1[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel1[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel1[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel1[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel1[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel1[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel1[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel1[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel1[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel1[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel1),
		.Data_Out(add_k1_Data_Out),
		.Valid_Out(add_kernel1_Valid_Out)
	);
	Batch_Norm bn_kernel1(
		.Data_A(32'b00111110100100001100000110001110),
		.Data_B(32'b00111110110010111111000010111011),
		.Data_In(add_k1_Data_Out),
		.Valid_In(add_kernel1_Valid_Out),
		.Data_Out(bn1_Data_Out),
		.Valid_Out(bn1_Valid_Out)
	);
	Relu_Core rl_kernel1(
		.Data_In(bn1_Data_Out),
		.Valid_In(bn1_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT-1:0]),
		.Valid_Out(rl1_Valid_Out)
	);
//////////KERNEL2//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111111000010101110110001000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111110101011111100001000101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110111010110110010100101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110100001110010010001000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111101100110001111000110110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110100101010000100000000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111110111010101011110011001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111110101111111011101110110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111100001111010001100000010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111100011100001110010000100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111101111011111100000111110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111100101110010100100110011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110100000101110001011101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111110101110100001110100111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110100111101010011010101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111110110110100011110111111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111101011100010110100010000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110011101110000110110000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110111101000111011111111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111111001100101110110001100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110101000110100001100101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111110101101000001010000110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111110110000001011110101110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111110111000001100101100000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111110010001001111001100000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111111001011110110011100010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110111100010010111000101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111100110100010100010100110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111110000100011010001111100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110100000001111101001001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111110100001010001001001001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111111010001000000100110000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel2_Valid_Out)
	);
	Adder_32input add_k2(
		.Data1(Data_Out_Kernel2[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel2[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel2[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel2[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel2[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel2[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel2[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel2[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel2[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel2[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel2[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel2[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel2[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel2[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel2[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel2[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel2[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel2[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel2[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel2[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel2[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel2[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel2[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel2[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel2[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel2[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel2[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel2[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel2[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel2[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel2[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel2[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel2),
		.Data_Out(add_k2_Data_Out),
		.Valid_Out(add_kernel2_Valid_Out)
	);
	Batch_Norm bn_kernel2(
		.Data_A(32'b00111110100000000111110100000001),
		.Data_B(32'b00111111100101011101111001111110),
		.Data_In(add_k2_Data_Out),
		.Valid_In(add_kernel2_Valid_Out),
		.Data_Out(bn2_Data_Out),
		.Valid_Out(bn2_Valid_Out)
	);
	Relu_Core rl_kernel2(
		.Data_In(bn2_Data_Out),
		.Valid_In(bn2_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Valid_Out(rl2_Valid_Out)
	);
//////////KERNEL3//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111110110010000011110101011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111101000011110100101101111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110101100010100111001010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111100110010000110011010100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111110010110011101110100100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111110100010110111000000001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111110100001110111000010001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111100110100100100110110011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111011100111011101111010001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110010010011110010000100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111111000010001100001100011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110110110100100011011101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110100000010001101000100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111100111111111001001000101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110001000110111011111011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111110110110100001011000010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110010010110101000111101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111111000110001011000110010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110001101100001100100101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110001101111000001000110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110000010001000111110110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111110111110001001011010110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111110001101011111000111111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111110011000011110010100101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111110001100010101000111000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111110011110100011111000010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111111001101010101100111110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111111000101010101100100000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111110111111011011101110100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110011011100110011111110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111111001111110011100111110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111110011111001101001000010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel3_Valid_Out)
	);
	Adder_32input add_k3(
		.Data1(Data_Out_Kernel3[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel3[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel3[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel3[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel3[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel3[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel3[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel3[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel3[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel3[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel3[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel3[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel3[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel3[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel3[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel3[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel3[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel3[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel3[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel3[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel3[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel3[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel3[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel3[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel3[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel3[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel3[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel3[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel3[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel3[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel3[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel3[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel3),
		.Data_Out(add_k3_Data_Out),
		.Valid_Out(add_kernel3_Valid_Out)
	);
	Batch_Norm bn_kernel3(
		.Data_A(32'b00111110010101110101110000110010),
		.Data_B(32'b00111110110010011001100010111001),
		.Data_In(add_k3_Data_Out),
		.Valid_In(add_kernel3_Valid_Out),
		.Data_Out(bn3_Data_Out),
		.Valid_Out(bn3_Valid_Out)
	);
	Relu_Core rl_kernel3(
		.Data_In(bn3_Data_Out),
		.Valid_In(bn3_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(rl3_Valid_Out)
	);
//////////KERNEL4//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110000001110010000000001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110011100110000110110100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111101011100000001001010100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111100111010000000001010110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111111001000110000101001110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110011101100000100101001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111110110001100110100100100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111111000111001111001011011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110111000000000100011010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111111000000001100011000100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110110001100010101010010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111101110100101111001000000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111110000111101101110000011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111110011011001101011000010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111111000100111001100000101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111100010110000011101010001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111111000010110101001111100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110011011111100000110010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111110011001111000000110110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111110011100100010111001010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110110000101101110001010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111110000110001010111110111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110010111111011101001111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111110000011100001011000000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111110100001110110110011001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110100110101000111110101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111111000100101100100011010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111111001001110010001101111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111110110111011110011000111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111101110000011111100110011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111110001001010110010100011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111111010111001101111101110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel4_Valid_Out)
	);
	Adder_32input add_k4(
		.Data1(Data_Out_Kernel4[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel4[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel4[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel4[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel4[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel4[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel4[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel4[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel4[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel4[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel4[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel4[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel4[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel4[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel4[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel4[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel4[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel4[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel4[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel4[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel4[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel4[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel4[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel4[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel4[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel4[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel4[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel4[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel4[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel4[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel4[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel4[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel4),
		.Data_Out(add_k4_Data_Out),
		.Valid_Out(add_kernel4_Valid_Out)
	);
	Batch_Norm bn_kernel4(
		.Data_A(32'b00111110100110011110001110100010),
		.Data_B(32'b00111111100111111011101011000011),
		.Data_In(add_k4_Data_Out),
		.Valid_In(add_kernel4_Valid_Out),
		.Data_Out(bn4_Data_Out),
		.Valid_Out(bn4_Valid_Out)
	);
	Relu_Core rl_kernel4(
		.Data_In(bn4_Data_Out),
		.Valid_In(bn4_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(rl4_Valid_Out)
	);
//////////KERNEL5//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110011111000000011011101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111110101010110011010101011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110110000100010011000011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111111001000111100100000100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111101101001000000011000000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111101011000111011111010010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111101110001111000111100100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111110100111101101011001110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110101010101100000111010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111101001101000010100010111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110101001110100010111100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111101101110000110100101110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111111010000000000011110101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111110011110101101100101100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111101111001001110111100111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111111000101010100001101010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111101000100001001001111101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111110000100110011100001111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111000000010110110110110110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111110000011010000000101000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110110101101101110110101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111110000001001011111111010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110100111111001100100100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111110001011100011101101100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111111001011011100100010110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111111011001111110011110010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111110010110011100110111011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110000100010010010010111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111111000100011001111001000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111111001100011000011111000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111110000100111101100001001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111011101001011010101110011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel5_Valid_Out)
	);
	Adder_32input add_k5(
		.Data1(Data_Out_Kernel5[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel5[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel5[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel5[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel5[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel5[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel5[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel5[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel5[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel5[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel5[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel5[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel5[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel5[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel5[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel5[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel5[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel5[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel5[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel5[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel5[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel5[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel5[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel5[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel5[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel5[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel5[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel5[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel5[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel5[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel5[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel5[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel5),
		.Data_Out(add_k5_Data_Out),
		.Valid_Out(add_kernel5_Valid_Out)
	);
	Batch_Norm bn_kernel5(
		.Data_A(32'b00111110100100000110110100010110),
		.Data_B(32'b10111110110000111101000100111000),
		.Data_In(add_k5_Data_Out),
		.Valid_In(add_kernel5_Valid_Out),
		.Data_Out(bn5_Data_Out),
		.Valid_Out(bn5_Valid_Out)
	);
	Relu_Core rl_kernel5(
		.Data_In(bn5_Data_Out),
		.Valid_In(bn5_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(rl5_Valid_Out)
	);
//////////KERNEL6//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111111000110000011000010011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111110101110111010001010010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111111001011001010101001110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111101110011000011001011011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111101010000110100011001100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110000101101001011111100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111111010000110101000110011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111110100111111101011001011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111101110101010110000011100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111111000000100010000010100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111101111010110011010000101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110011001011110011010000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111110000010100100110101101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111101101001010110011001101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110111101011000000101010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111111000101010010010100101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111110100111010011000111111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110111011011000001101111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110110011100011011100000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111110000100100000101101011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111101110101110011000000000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111110110001000100011110010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110001111111000010110101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111111010001100001000010010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111110110011111100111011001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110100010001001110100100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111110100000000101111001111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111101100101110001110111111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111110000000101101011000011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111110101011010101001110000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111110011011010000011010011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111110010011111110101011001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel6_Valid_Out)
	);
	Adder_32input add_k6(
		.Data1(Data_Out_Kernel6[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel6[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel6[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel6[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel6[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel6[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel6[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel6[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel6[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel6[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel6[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel6[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel6[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel6[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel6[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel6[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel6[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel6[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel6[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel6[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel6[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel6[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel6[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel6[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel6[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel6[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel6[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel6[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel6[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel6[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel6[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel6[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel6),
		.Data_Out(add_k6_Data_Out),
		.Valid_Out(add_kernel6_Valid_Out)
	);
	Batch_Norm bn_kernel6(
		.Data_A(32'b00111110101000000001001010011011),
		.Data_B(32'b00111110100111111000100000001000),
		.Data_In(add_k6_Data_Out),
		.Valid_In(add_kernel6_Valid_Out),
		.Data_Out(bn6_Data_Out),
		.Valid_Out(bn6_Valid_Out)
	);
	Relu_Core rl_kernel6(
		.Data_In(bn6_Data_Out),
		.Valid_In(bn6_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(rl6_Valid_Out)
	);
//////////KERNEL7//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110010001011110000011110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110101100011101000011000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110010001101000101110110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110101010000011110000001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111110010100001011001011010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111101110101011001111101111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111110110000001001000100000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111110100110110110000111101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111110101011001001010100010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111111000111001100000010001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111110010010101110101100101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111101110110011001000110100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111111000010010000110010101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111110101001010110100000110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111101111100010001101011101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111110010110111100100010000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111110100100111101000111000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110010010100010110101101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110001101110100001101101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111110011100001111111101111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111101110001100001000110110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111111001011111111110110100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111101000111000010011010100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111101101100000110001001000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111110011110000100110001000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111110100101010010010000111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111110100110111001110001010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111100101100001000100101110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111111001010000100101101010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110010010111111001000111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111111011111100100111101000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110101111001001010010101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel7_Valid_Out)
	);
	Adder_32input add_k7(
		.Data1(Data_Out_Kernel7[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel7[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel7[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel7[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel7[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel7[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel7[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel7[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel7[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel7[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel7[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel7[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel7[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel7[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel7[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel7[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel7[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel7[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel7[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel7[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel7[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel7[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel7[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel7[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel7[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel7[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel7[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel7[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel7[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel7[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel7[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel7[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel7),
		.Data_Out(add_k7_Data_Out),
		.Valid_Out(add_kernel7_Valid_Out)
	);
	Batch_Norm bn_kernel7(
		.Data_A(32'b00111110010110110110000010010001),
		.Data_B(32'b00111111001110000101110110101011),
		.Data_In(add_k7_Data_Out),
		.Valid_In(add_kernel7_Valid_Out),
		.Data_Out(bn7_Data_Out),
		.Valid_Out(bn7_Valid_Out)
	);
	Relu_Core rl_kernel7(
		.Data_In(bn7_Data_Out),
		.Valid_In(bn7_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(rl7_Valid_Out)
	);
//////////KERNEL8//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111110101111001000010101011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111101100101000100110010111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110000010101110011101011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111101101100001000001110000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111100110110111101011000010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111101010010111001100001101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111110011010000010101101101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111110010110000011011101010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111101010010011110101110101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111110101011101110011011101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111110001010111111001010111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111111001100001101001111100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111110110111111000111010110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111110001111001001100101100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111111000110011100100010111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111110100001111110001110110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110101011010010100010011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110011111000100001110101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111101111110100101001100000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111111000001000011100001001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111011100010000110011010010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111110010010000111001100101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111110101111001011100001111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111111100011000100100111001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111110011101101000110010110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111101000010111111100010100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110100110111001000011110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111111000110001000011101001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111111010010001000100101000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110001100101010100001011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111110000101101000111110111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111100001111011001111010010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel8_Valid_Out)
	);
	Adder_32input add_k8(
		.Data1(Data_Out_Kernel8[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel8[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel8[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel8[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel8[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel8[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel8[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel8[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel8[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel8[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel8[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel8[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel8[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel8[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel8[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel8[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel8[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel8[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel8[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel8[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel8[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel8[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel8[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel8[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel8[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel8[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel8[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel8[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel8[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel8[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel8[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel8[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel8),
		.Data_Out(add_k8_Data_Out),
		.Valid_Out(add_kernel8_Valid_Out)
	);
	Batch_Norm bn_kernel8(
		.Data_A(32'b00111110011001011101111111110011),
		.Data_B(32'b00111110111111101100101100110001),
		.Data_In(add_k8_Data_Out),
		.Valid_In(add_kernel8_Valid_Out),
		.Data_Out(bn8_Data_Out),
		.Valid_Out(bn8_Valid_Out)
	);
	Relu_Core rl_kernel8(
		.Data_In(bn8_Data_Out),
		.Valid_In(bn8_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(rl8_Valid_Out)
	);
//////////KERNEL9//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111110111001110011101111101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110001011110101101110011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110010000001111010011111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111011100000010010001101110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111110111111001011100110011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111100011001111101000110011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111101110110111111100100110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111110010011011111110100010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111101000011000110101110110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110100110000111111010001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111100110110010010100101000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111101110110111100110100100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111111100001111011010110110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111110110000000000111110100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110111110010010101110011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111110010000100101010000100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110101100110100111100011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111110101011001011101110001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110100110110100100000000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111100110100110010000111110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111111001101011000101101111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111101000000111001001110011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111111001001110010110111001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111111000001000100011111100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111110110000110100111100110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111101010111001000000101110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111100001110011100011111110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111110011011100110110001010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111110110000111000011000100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111110111110111000100001110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111110110011001010100011011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110011000011111100110101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel9_Valid_Out)
	);
	Adder_32input add_k9(
		.Data1(Data_Out_Kernel9[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel9[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel9[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel9[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel9[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel9[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel9[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel9[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel9[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel9[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel9[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel9[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel9[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel9[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel9[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel9[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel9[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel9[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel9[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel9[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel9[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel9[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel9[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel9[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel9[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel9[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel9[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel9[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel9[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel9[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel9[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel9[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel9),
		.Data_Out(add_k9_Data_Out),
		.Valid_Out(add_kernel9_Valid_Out)
	);
	Batch_Norm bn_kernel9(
		.Data_A(32'b00111110101110000111111101101100),
		.Data_B(32'b10111110010101110011000011010101),
		.Data_In(add_k9_Data_Out),
		.Valid_In(add_kernel9_Valid_Out),
		.Data_Out(bn9_Data_Out),
		.Valid_Out(bn9_Valid_Out)
	);
	Relu_Core rl_kernel9(
		.Data_In(bn9_Data_Out),
		.Valid_In(bn9_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(rl9_Valid_Out)
	);
//////////KERNEL10//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111101101101010010100100010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111110010000001011001101100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110111000000000001101101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111101000000101111001100110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111110000100010000110000001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111110110101101111000111100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111110101000100101011111100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111111100000101110110101111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111110100110011001011111110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111101111000010100101101011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111111000011101101000100100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110110011110010101000011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111110101101001110001101001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111101001110101111101110001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111101101000001010101001001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111100111101110000010011100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110101000011110000000000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110011110100100000100011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111110010110100010111001110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111111010001101010001100110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110001000111110100101101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111110111100111010111111011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110100100011100011111000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111110010100010000000000001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111110100010110000100010001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111100101111001111001010110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110010100101000110001000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111111010101010010001010100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111110001000001010100000010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111101000011001110011011000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111101000110110001010110101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111110101000011001010010010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel10_Valid_Out)
	);
	Adder_32input add_k10(
		.Data1(Data_Out_Kernel10[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel10[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel10[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel10[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel10[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel10[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel10[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel10[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel10[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel10[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel10[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel10[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel10[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel10[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel10[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel10[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel10[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel10[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel10[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel10[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel10[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel10[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel10[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel10[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel10[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel10[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel10[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel10[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel10[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel10[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel10[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel10[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel10),
		.Data_Out(add_k10_Data_Out),
		.Valid_Out(add_kernel10_Valid_Out)
	);
	Batch_Norm bn_kernel10(
		.Data_A(32'b00111110100100100010010101010111),
		.Data_B(32'b00111110000011010011101110110001),
		.Data_In(add_k10_Data_Out),
		.Valid_In(add_kernel10_Valid_Out),
		.Data_Out(bn10_Data_Out),
		.Valid_Out(bn10_Valid_Out)
	);
	Relu_Core rl_kernel10(
		.Data_In(bn10_Data_Out),
		.Valid_In(bn10_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(rl10_Valid_Out)
	);
//////////KERNEL11//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111110100110011001001111011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111101001100010111011110110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110000010101011010101110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111100100100111011110010110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111110001100001100110100001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111101110011111101010101011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111110001110111101010001101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111111001001001000110100011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111111010011100111110001110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111111000111111000010011010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111111100100000010011110110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110100111100101011101000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111101100101100100100011100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111110000110111110000110111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110101011011110100001010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111110101000010100010011111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111101101111001100111111001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111110011010100111100010110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110100000000000111101000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111101111101010010110011011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110101111110111111110011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111110001011001011010000010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111110101011101111100011111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111101100100111011101010010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111110111000110110000110010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110101001011001000001010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111011110110100100001100101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111111001110010000110001010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111101101101001000111011000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110011000000011101111100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111110100111111011110100111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111101101010101010010111101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel11_Valid_Out)
	);
	Adder_32input add_k11(
		.Data1(Data_Out_Kernel11[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel11[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel11[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel11[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel11[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel11[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel11[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel11[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel11[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel11[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel11[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel11[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel11[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel11[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel11[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel11[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel11[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel11[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel11[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel11[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel11[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel11[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel11[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel11[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel11[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel11[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel11[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel11[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel11[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel11[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel11[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel11[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel11),
		.Data_Out(add_k11_Data_Out),
		.Valid_Out(add_kernel11_Valid_Out)
	);
	Batch_Norm bn_kernel11(
		.Data_A(32'b00111110100101011010110110000110),
		.Data_B(32'b00111111100000101100100110101001),
		.Data_In(add_k11_Data_Out),
		.Valid_In(add_kernel11_Valid_Out),
		.Data_Out(bn11_Data_Out),
		.Valid_Out(bn11_Valid_Out)
	);
	Relu_Core rl_kernel11(
		.Data_In(bn11_Data_Out),
		.Valid_In(bn11_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(rl11_Valid_Out)
	);
//////////KERNEL12//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111111001001111010110011011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111110111001011101111011011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111101100111010001110000101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110010101110010110110001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111110101011101000000111000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111110001111000001110000111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111110101000010001001100101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111110100011010111111101001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111111000100011101010111111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111111001110010110101111000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110100000001101111110111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111110101001001100001010001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111110100111010110101010101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111111000001100111110111011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110101011001010010000000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111101111011011100010100111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111111000001011110100100000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111110000000001011100011000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111110001001011110011110011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111101101100110011000000110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111101111001000000110101101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111100001110000011000011001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111111001100001111100001110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111011110011111010001011101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111110010011011001111000010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111110101100011100011000111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111110001100111000111010111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110111010010001010100101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111110111000100011101001001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110100111111111100111111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111101111111101001010100010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110000100100000101000101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel12_Valid_Out)
	);
	Adder_32input add_k12(
		.Data1(Data_Out_Kernel12[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel12[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel12[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel12[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel12[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel12[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel12[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel12[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel12[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel12[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel12[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel12[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel12[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel12[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel12[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel12[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel12[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel12[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel12[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel12[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel12[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel12[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel12[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel12[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel12[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel12[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel12[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel12[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel12[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel12[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel12[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel12[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel12),
		.Data_Out(add_k12_Data_Out),
		.Valid_Out(add_kernel12_Valid_Out)
	);
	Batch_Norm bn_kernel12(
		.Data_A(32'b00111110111000110011101101101111),
		.Data_B(32'b10111110010101011100100001110110),
		.Data_In(add_k12_Data_Out),
		.Valid_In(add_kernel12_Valid_Out),
		.Data_Out(bn12_Data_Out),
		.Valid_Out(bn12_Valid_Out)
	);
	Relu_Core rl_kernel12(
		.Data_In(bn12_Data_Out),
		.Valid_In(bn12_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(rl12_Valid_Out)
	);
//////////KERNEL13//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111110101110100101110001000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111101001010110011110010111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110011100010001010001010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110100001001111000101101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111111001001110011011100010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111101011001011010110100101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111111000100010001111101010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111101110111110011111110001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111001010011000111101000101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110101100011110101111001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111101111001011111100101101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111111000101010001011110001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111111011100101010100010101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111110000100100100101000101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111101111101011101101000011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111110100000001001110101110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110110011010111001110010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111110100111100111110001110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111110001001011011011010111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111110010010001000100101011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110011101000100011111011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111110000000100101011110111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110000100100101000101001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111111000101111110110111100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111110011011111100010010001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111100110000111111111110100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111111000101010011111111111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111110001101010110000010010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111111001000010000000001001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111100100110100010101010111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111101100110010011010111110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110101001101011111100101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel13_Valid_Out)
	);
	Adder_32input add_k13(
		.Data1(Data_Out_Kernel13[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel13[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel13[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel13[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel13[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel13[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel13[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel13[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel13[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel13[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel13[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel13[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel13[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel13[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel13[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel13[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel13[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel13[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel13[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel13[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel13[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel13[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel13[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel13[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel13[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel13[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel13[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel13[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel13[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel13[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel13[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel13[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel13),
		.Data_Out(add_k13_Data_Out),
		.Valid_Out(add_kernel13_Valid_Out)
	);
	Batch_Norm bn_kernel13(
		.Data_A(32'b00111110100010100010100010010000),
		.Data_B(32'b00111101100000110111001000011001),
		.Data_In(add_k13_Data_Out),
		.Valid_In(add_kernel13_Valid_Out),
		.Data_Out(bn13_Data_Out),
		.Valid_Out(bn13_Valid_Out)
	);
	Relu_Core rl_kernel13(
		.Data_In(bn13_Data_Out),
		.Valid_In(bn13_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(rl13_Valid_Out)
	);
//////////KERNEL14//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111110000010101111100001010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111110000000101000111110110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110100011101011101110001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111111000010100100100111011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111110101000110010100010010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111100101101111111101101110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111111000011001101101110101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111111000110000000110100101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111111001110010001100001101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111101011011100011111111100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111110000001101100011111101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110000000001001111111011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111110001000011101011101111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111101010111101001100010000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110101000011101011111100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111110100010101000100010110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111010110010010110010100111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111101110111100000011111010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111111100000100001110110010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111111001000011001000001111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110000011010011000100111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111101111100101001111000001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110110001111101000011100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111101101111011111110100000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111100000100010011001111111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111100100110010001011000000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111101111101011001101111001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111101001111111010101000101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111111010000111011011110010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111101101011111011010100111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111110110001100101101010000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111100101100011100101001001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel14_Valid_Out)
	);
	Adder_32input add_k14(
		.Data1(Data_Out_Kernel14[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel14[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel14[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel14[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel14[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel14[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel14[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel14[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel14[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel14[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel14[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel14[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel14[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel14[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel14[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel14[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel14[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel14[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel14[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel14[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel14[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel14[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel14[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel14[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel14[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel14[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel14[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel14[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel14[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel14[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel14[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel14[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel14),
		.Data_Out(add_k14_Data_Out),
		.Valid_Out(add_kernel14_Valid_Out)
	);
	Batch_Norm bn_kernel14(
		.Data_A(32'b00111110100001111111110100111110),
		.Data_B(32'b00111111001001110100001111101001),
		.Data_In(add_k14_Data_Out),
		.Valid_In(add_kernel14_Valid_Out),
		.Data_Out(bn14_Data_Out),
		.Valid_Out(bn14_Valid_Out)
	);
	Relu_Core rl_kernel14(
		.Data_In(bn14_Data_Out),
		.Valid_In(bn14_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(rl14_Valid_Out)
	);
//////////KERNEL15//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110000100010011111110000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111101111000101100100101111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111101111010010001101001001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111111000101100001101111001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111110011001001111111011101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111110100101010000101010101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111101110100101111101011101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111111010011100111011110011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110100011100001010111100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111101110101111011100101110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110101000111001101100110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111101111110110001100110110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111100110110111111011101011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111110101001011101110010110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110101010011111001100111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111111000110011000010110110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111110101010111011010011000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111111000110101011000011000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110111100100011111010011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110100010001100100111010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110101111011101011001011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111110000011000011101101111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111101110010100110100110110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111111001110011110000011111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111101000000010010011001000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111110010010100110101000000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111111001100111111110000110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110011100100000100111011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111101111100010100101011110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111110000110010011011000111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111110111001011110100101101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111101011100110100111110010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel15_Valid_Out)
	);
	Adder_32input add_k15(
		.Data1(Data_Out_Kernel15[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel15[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel15[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel15[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel15[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel15[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel15[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel15[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel15[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel15[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel15[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel15[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel15[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel15[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel15[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel15[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel15[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel15[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel15[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel15[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel15[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel15[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel15[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel15[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel15[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel15[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel15[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel15[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel15[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel15[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel15[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel15[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel15),
		.Data_Out(add_k15_Data_Out),
		.Valid_Out(add_kernel15_Valid_Out)
	);
	Batch_Norm bn_kernel15(
		.Data_A(32'b00111110110001010110100011001111),
		.Data_B(32'b00111111110100110100101011111001),
		.Data_In(add_k15_Data_Out),
		.Valid_In(add_kernel15_Valid_Out),
		.Data_Out(bn15_Data_Out),
		.Valid_Out(bn15_Valid_Out)
	);
	Relu_Core rl_kernel15(
		.Data_In(bn15_Data_Out),
		.Valid_In(bn15_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(rl15_Valid_Out)
	);
//////////KERNEL16//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111111010110101001111101010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110010000100100100001011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110010111011111010010100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111101101111100001101001011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111100110101001001110101011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111111000000000011001011111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111101101100011111100110111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111111000111111101001000110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111101110010010111111110111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110111010111010101100100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110011000001110110010111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111110111001000000111101000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111111010110101010101110111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111101100111010101010110010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111101000100101100001101100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111111001010010000110011010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111110101011111010111100011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110100011110101011101111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110000001100000010011011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111110011110000000110001100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111101110011010010000000111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111110011000111110100000001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110000101100110011111110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111100111011010110110011001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111110011100100011111100011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111101101100000100011011110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110100011100101000010111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111111001110101100001101000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111101111111110100000101100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111101101000000000011111111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111110011111111101010111010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111111000101001111101010101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel16_Valid_Out)
	);
	Adder_32input add_k16(
		.Data1(Data_Out_Kernel16[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel16[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel16[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel16[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel16[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel16[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel16[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel16[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel16[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel16[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel16[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel16[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel16[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel16[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel16[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel16[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel16[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel16[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel16[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel16[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel16[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel16[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel16[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel16[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel16[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel16[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel16[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel16[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel16[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel16[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel16[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel16[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel16),
		.Data_Out(add_k16_Data_Out),
		.Valid_Out(add_kernel16_Valid_Out)
	);
	Batch_Norm bn_kernel16(
		.Data_A(32'b00111110100010111110000011010110),
		.Data_B(32'b00111111100101111100100011000101),
		.Data_In(add_k16_Data_Out),
		.Valid_In(add_kernel16_Valid_Out),
		.Data_Out(bn16_Data_Out),
		.Valid_Out(bn16_Valid_Out)
	);
	Relu_Core rl_kernel16(
		.Data_In(bn16_Data_Out),
		.Valid_In(bn16_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(rl16_Valid_Out)
	);
//////////KERNEL17//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111100001011011000111101001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110001101011101010101011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111101111100101110100000110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110001001001111101010111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111110100111011001001000101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111111000101110000000001101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111110001001000011001100111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111110111011111000010111101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110100111100100000000100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110111111000010010000101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110010110100110101111111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110100011010101101101011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110101011110011010011001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111101101001011110101010001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110100010111100111010011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111101110110101111011001100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111011001110011101001111010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110100001001010111000001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111111000111101111011011001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111110111100100000100111101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111111010100001001000001010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111110101100001111011110100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111101111000010010101000001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111111001010001010001001110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111111001000110011001110101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111101100011001010111011000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110000000110001111011111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111101100110001101001000100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111111000011000111100110010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111110101000110011101011100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111101101010100110000001110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111100100000111000111111000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel17_Valid_Out)
	);
	Adder_32input add_k17(
		.Data1(Data_Out_Kernel17[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel17[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel17[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel17[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel17[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel17[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel17[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel17[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel17[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel17[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel17[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel17[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel17[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel17[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel17[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel17[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel17[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel17[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel17[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel17[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel17[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel17[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel17[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel17[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel17[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel17[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel17[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel17[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel17[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel17[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel17[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel17[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel17),
		.Data_Out(add_k17_Data_Out),
		.Valid_Out(add_kernel17_Valid_Out)
	);
	Batch_Norm bn_kernel17(
		.Data_A(32'b00111110100100111000111111111001),
		.Data_B(32'b00111110101001010110001011000000),
		.Data_In(add_k17_Data_Out),
		.Valid_In(add_kernel17_Valid_Out),
		.Data_Out(bn17_Data_Out),
		.Valid_Out(bn17_Valid_Out)
	);
	Relu_Core rl_kernel17(
		.Data_In(bn17_Data_Out),
		.Valid_In(bn17_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(rl17_Valid_Out)
	);
//////////KERNEL18//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111110100110000011011010110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111111001000100001111000011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110110010011110111000111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111111001010100001001101011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111101100100100010111000010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111110001001101011000110001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111110001110111100010011100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111101111111111001100101000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110000010100001001010000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110110101101100111100111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111101101001110100010111001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110101100000001001001000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111101011001110010111110101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111110101110000001001010010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111111100101111000001000010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111111000100000000101000001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110110100100110111111000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111100010010100001001110110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111111001010010111111010110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111101011011010010000101000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110100100010011000001101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111110011000100101010100000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111101110100110111000001111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111101111001001100001100111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111110011111000000111100001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111110100011000011100101110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111111001011000001101100000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111110000000001011101110010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111110010001101000111110010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110000101001011011111110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111101111101110001111011111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110010011110100101011011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel18_Valid_Out)
	);
	Adder_32input add_k18(
		.Data1(Data_Out_Kernel18[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel18[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel18[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel18[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel18[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel18[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel18[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel18[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel18[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel18[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel18[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel18[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel18[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel18[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel18[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel18[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel18[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel18[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel18[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel18[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel18[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel18[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel18[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel18[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel18[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel18[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel18[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel18[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel18[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel18[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel18[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel18[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel18),
		.Data_Out(add_k18_Data_Out),
		.Valid_Out(add_kernel18_Valid_Out)
	);
	Batch_Norm bn_kernel18(
		.Data_A(32'b00111110010101100011001010010110),
		.Data_B(32'b00111101000010000101101101001010),
		.Data_In(add_k18_Data_Out),
		.Valid_In(add_kernel18_Valid_Out),
		.Data_Out(bn18_Data_Out),
		.Valid_Out(bn18_Valid_Out)
	);
	Relu_Core rl_kernel18(
		.Data_In(bn18_Data_Out),
		.Valid_In(bn18_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(rl18_Valid_Out)
	);
//////////KERNEL19//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111101101000011101100101110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111100011100011000101000100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110100001001010101110011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110100111011001111001110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111101101011101010000011010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110110000100111111010101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111100100110110011100011100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111110110110110000100010010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110110111100101100000101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110100010010001101111010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111111010001101111101010111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111111001000100110000000000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110011110111010010011111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111110011000010000110101010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110001001000100110001001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111110101011010011110001111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110000100111110110111110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111101101011111111000100011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111100110010110001111010001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111110000110101011100101110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110111111100101100001001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111111010010110011100011011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111110101001010010111110100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111110111000101001110000001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111110110101000101100000111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110000101001110111011110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110100011010110011011000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110110010110011111110011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111111010010101101010100110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111101101110111011010110011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111110010100001001011011001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111110100101110001010011110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel19_Valid_Out)
	);
	Adder_32input add_k19(
		.Data1(Data_Out_Kernel19[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel19[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel19[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel19[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel19[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel19[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel19[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel19[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel19[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel19[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel19[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel19[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel19[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel19[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel19[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel19[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel19[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel19[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel19[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel19[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel19[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel19[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel19[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel19[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel19[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel19[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel19[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel19[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel19[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel19[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel19[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel19[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel19),
		.Data_Out(add_k19_Data_Out),
		.Valid_Out(add_kernel19_Valid_Out)
	);
	Batch_Norm bn_kernel19(
		.Data_A(32'b00111110011101001011111110000100),
		.Data_B(32'b00111011101100111100000101000000),
		.Data_In(add_k19_Data_Out),
		.Valid_In(add_kernel19_Valid_Out),
		.Data_Out(bn19_Data_Out),
		.Valid_Out(bn19_Valid_Out)
	);
	Relu_Core rl_kernel19(
		.Data_In(bn19_Data_Out),
		.Valid_In(bn19_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(rl19_Valid_Out)
	);
//////////KERNEL20//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110110000100011111010001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111101001111011110111101110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111111011111100000110101111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110010010110100101101110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111100000001001101100111110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111101001100110101011111000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111110010011000110011110101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111101101110001100101010010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110101110001111010010011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110110010111111110101011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111111011000101101000100110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111101110111111110111100100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111101101001011001001011100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111100100001101110011010000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111111000100000001110010100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111101111010011101110010110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111111001001001101001111011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111110001001101111111011100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111110100100100111011110101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111100100011111011110101011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111111001011010010100000010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111101101100100001011001111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111111001011101001010100100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111101101000010111010111101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111110101001000011110010101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111110110100111100100001100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111100110110101000101100110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110100010000101101011010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111110001011010110000000100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111101111001101010110001011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111110101101110011100000111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110000011100111001010101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel20_Valid_Out)
	);
	Adder_32input add_k20(
		.Data1(Data_Out_Kernel20[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel20[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel20[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel20[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel20[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel20[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel20[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel20[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel20[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel20[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel20[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel20[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel20[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel20[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel20[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel20[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel20[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel20[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel20[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel20[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel20[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel20[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel20[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel20[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel20[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel20[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel20[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel20[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel20[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel20[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel20[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel20[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel20),
		.Data_Out(add_k20_Data_Out),
		.Valid_Out(add_kernel20_Valid_Out)
	);
	Batch_Norm bn_kernel20(
		.Data_A(32'b00111110011111010010010110110100),
		.Data_B(32'b00111110111100010010100010010101),
		.Data_In(add_k20_Data_Out),
		.Valid_In(add_kernel20_Valid_Out),
		.Data_Out(bn20_Data_Out),
		.Valid_Out(bn20_Valid_Out)
	);
	Relu_Core rl_kernel20(
		.Data_In(bn20_Data_Out),
		.Valid_In(bn20_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(rl20_Valid_Out)
	);
//////////KERNEL21//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111110100010001000000011000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110010000000110001111001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110101110101010001110100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111100011011101011000001110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111110101000000001011100111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111100100101000000111000110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111110000001111001010101110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111111010111011010011011011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111110010101001011001001111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110110001100000100101000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111101100010000001101111111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110110011111010100010101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110010100010110000110011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111101001110001101111111011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110110010110100011111100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111110001110111100111000100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111101101000110110011100001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111111000100001101110111000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111111000110111110111000000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110100101000000111001000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110010001101000111110001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111111000110000100100100110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110010010010111000110100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111110001100100110110100101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111110110001111001001101010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111110001101010110011000101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111110100101100000000110111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111110010101110000010001111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111110000110110001110001011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111110001100000111100110100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111111010111010011110101011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111101001110001100011110010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel21_Valid_Out)
	);
	Adder_32input add_k21(
		.Data1(Data_Out_Kernel21[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel21[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel21[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel21[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel21[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel21[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel21[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel21[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel21[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel21[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel21[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel21[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel21[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel21[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel21[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel21[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel21[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel21[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel21[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel21[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel21[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel21[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel21[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel21[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel21[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel21[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel21[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel21[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel21[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel21[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel21[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel21[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel21),
		.Data_Out(add_k21_Data_Out),
		.Valid_Out(add_kernel21_Valid_Out)
	);
	Batch_Norm bn_kernel21(
		.Data_A(32'b00111110011100110111101011011010),
		.Data_B(32'b00111101000011001011110111010111),
		.Data_In(add_k21_Data_Out),
		.Valid_In(add_kernel21_Valid_Out),
		.Data_Out(bn21_Data_Out),
		.Valid_Out(bn21_Valid_Out)
	);
	Relu_Core rl_kernel21(
		.Data_In(bn21_Data_Out),
		.Valid_In(bn21_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(rl21_Valid_Out)
	);
//////////KERNEL22//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111111001100110000111110110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111111010001110110100100111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111101100101011000011111101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111101101100010101001001011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111110100010011001000010110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110001111110010011110001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111111001001011101111101111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111100010110111101110000000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111111000110010110111001010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110001101011011111011100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110001001100111110100011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111100111000001011011101101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110010010011000001111000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111111001011101101110011000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111010100100101000000011000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111110001101111001000010101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111101110010000000000101011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111100110000000010100101001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111111001000111111101010111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111101100100101000000000100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110110110100000000000110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111110110001110010001011011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110101101110111000010100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111110010101000000000000110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111101000010000000110111011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111111010001010010101011111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110100101001101111000001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111110000100110100001011011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111110010001110010110010000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110001010000101111010100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111110111010110000111110010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111101110010011011101111010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel22_Valid_Out)
	);
	Adder_32input add_k22(
		.Data1(Data_Out_Kernel22[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel22[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel22[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel22[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel22[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel22[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel22[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel22[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel22[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel22[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel22[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel22[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel22[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel22[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel22[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel22[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel22[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel22[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel22[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel22[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel22[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel22[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel22[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel22[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel22[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel22[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel22[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel22[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel22[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel22[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel22[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel22[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel22),
		.Data_Out(add_k22_Data_Out),
		.Valid_Out(add_kernel22_Valid_Out)
	);
	Batch_Norm bn_kernel22(
		.Data_A(32'b00111110010110100100110101100111),
		.Data_B(32'b00111101000001010110001001000100),
		.Data_In(add_k22_Data_Out),
		.Valid_In(add_kernel22_Valid_Out),
		.Data_Out(bn22_Data_Out),
		.Valid_Out(bn22_Valid_Out)
	);
	Relu_Core rl_kernel22(
		.Data_In(bn22_Data_Out),
		.Valid_In(bn22_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(rl22_Valid_Out)
	);
//////////KERNEL23//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110100010011000111010100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110111000001110111110100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111111000000100101100001100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111111000011100101111101101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111100100010111110001111100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111111000101001100001111010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111100001110011000001001000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111101010101000010101111000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110110000100101000100000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111101011010000011100001110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111101110101001000011100111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111101111010101011000111010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110111010110111001001011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111001100100010100101100001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110101101001010011111111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111110101000110011000101100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111110100010010101100001011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110110111000110111110001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111110101011010010000011011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110110010011001110111000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110110000110100101101110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111101110101001110101100011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110110111100100111100111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111110101100010011111000011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111110110000100110110010100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111101010101101101011010111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110100111011111001100101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111110100000011101000000001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111110100010100111000001010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111111010010010101110110010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111110101000111100100101100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111111001001101110101110111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel23_Valid_Out)
	);
	Adder_32input add_k23(
		.Data1(Data_Out_Kernel23[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel23[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel23[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel23[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel23[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel23[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel23[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel23[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel23[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel23[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel23[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel23[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel23[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel23[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel23[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel23[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel23[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel23[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel23[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel23[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel23[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel23[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel23[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel23[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel23[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel23[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel23[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel23[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel23[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel23[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel23[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel23[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel23),
		.Data_Out(add_k23_Data_Out),
		.Valid_Out(add_kernel23_Valid_Out)
	);
	Batch_Norm bn_kernel23(
		.Data_A(32'b00111110101001000000010100101110),
		.Data_B(32'b00111110100001101011110010111111),
		.Data_In(add_k23_Data_Out),
		.Valid_In(add_kernel23_Valid_Out),
		.Data_Out(bn23_Data_Out),
		.Valid_Out(bn23_Valid_Out)
	);
	Relu_Core rl_kernel23(
		.Data_In(bn23_Data_Out),
		.Valid_In(bn23_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(rl23_Valid_Out)
	);
//////////KERNEL24//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111110111110000001100111001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111110010100100011111011011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110001110100110010110011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110111011010010101100101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111110001111000011100110010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110101010111101111101011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111011111000100101101001010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111101101011100101000011000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110100111111101010101100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111110100000101010101110011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110100000111001011111111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111101000001010110110100010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111101111101110111000110111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111100110000101000010011110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110000000110111010001011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111110010000001001011001101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111101010111100101110110001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111111000011011001100110100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110111000000111001101010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111110011111110000101011011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111111001000110000000001011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111110000001011001100111110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111111000000100100110011011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111110010101101111101101001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111101111011010010111001101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110100111010011010000100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111111011011011111000011111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110101100010101000110111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111110101110000010000101000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110010010100011011100000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111100011000000101110000100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111111011001110101011010011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel24_Valid_Out)
	);
	Adder_32input add_k24(
		.Data1(Data_Out_Kernel24[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel24[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel24[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel24[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel24[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel24[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel24[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel24[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel24[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel24[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel24[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel24[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel24[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel24[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel24[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel24[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel24[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel24[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel24[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel24[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel24[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel24[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel24[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel24[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel24[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel24[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel24[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel24[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel24[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel24[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel24[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel24[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel24),
		.Data_Out(add_k24_Data_Out),
		.Valid_Out(add_kernel24_Valid_Out)
	);
	Batch_Norm bn_kernel24(
		.Data_A(32'b00111110101100000000100001011001),
		.Data_B(32'b00111110111101011010111100001101),
		.Data_In(add_k24_Data_Out),
		.Valid_In(add_kernel24_Valid_Out),
		.Data_Out(bn24_Data_Out),
		.Valid_Out(bn24_Valid_Out)
	);
	Relu_Core rl_kernel24(
		.Data_In(bn24_Data_Out),
		.Valid_In(bn24_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(rl24_Valid_Out)
	);
//////////KERNEL25//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110101101110010010001010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111110101001000110111010010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110011100101101011011000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111111000110000011111111010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111110100110110110010000001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111110011011001000001110101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111011100011010001100010001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111111000001011111101101000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110101110100111110010001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111101100000111100111010001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111110110100001101100100110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110110001110100100001011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111101100000000110100001110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111101110100111111100100101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110100010111100000001000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111101110100101000010011010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111101100111101111010110111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111110100000011010110101011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110010100000010111100100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110111110100010110000101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110000100100000011101100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111111010010111001111011111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110100101110000101110111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111110101010001010010101111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111101101011101010000011100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111101101111100110001011110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111101011111101101010111001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111110000101001000101101100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111110011000000010001101000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110100100111010000000010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111111011100001000001000100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111111000001110111001101110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel25_Valid_Out)
	);
	Adder_32input add_k25(
		.Data1(Data_Out_Kernel25[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel25[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel25[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel25[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel25[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel25[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel25[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel25[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel25[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel25[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel25[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel25[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel25[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel25[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel25[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel25[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel25[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel25[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel25[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel25[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel25[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel25[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel25[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel25[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel25[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel25[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel25[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel25[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel25[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel25[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel25[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel25[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel25),
		.Data_Out(add_k25_Data_Out),
		.Valid_Out(add_kernel25_Valid_Out)
	);
	Batch_Norm bn_kernel25(
		.Data_A(32'b00111110100100101101111000101110),
		.Data_B(32'b00111110010101111111100010110101),
		.Data_In(add_k25_Data_Out),
		.Valid_In(add_kernel25_Valid_Out),
		.Data_Out(bn25_Data_Out),
		.Valid_Out(bn25_Valid_Out)
	);
	Relu_Core rl_kernel25(
		.Data_In(bn25_Data_Out),
		.Valid_In(bn25_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(rl25_Valid_Out)
	);
//////////KERNEL26//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111110000001001011100101100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111111000011100111100101001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110111100011110011111101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111100100111000011000011000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111011111011011001011101100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111110010010110111011111001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111101110000011010111110010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111100000100000101011010010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111110101101011001110100100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111110100111100010011010110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111100000001111010001101111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110001100011000011001110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111101100110000110100011011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111110011101111111110011010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110000011100001111100100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111111000111010101110011110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111111000101111110101010001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111110001010110010000100111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111111000111010111110000001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111111000001001000110011001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110111011110111100111010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111110111100011100111011111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111011100110000011110101010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111110100001111101011001011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111110100011000111100100011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111110100101000010010100101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110011101010001110011011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110110011010101011110010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111111001000000110001010011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111110000000100001000101001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111110111000101001010111001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110110100010001011101001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel26_Valid_Out)
	);
	Adder_32input add_k26(
		.Data1(Data_Out_Kernel26[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel26[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel26[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel26[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel26[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel26[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel26[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel26[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel26[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel26[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel26[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel26[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel26[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel26[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel26[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel26[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel26[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel26[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel26[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel26[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel26[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel26[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel26[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel26[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel26[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel26[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel26[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel26[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel26[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel26[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel26[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel26[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel26),
		.Data_Out(add_k26_Data_Out),
		.Valid_Out(add_kernel26_Valid_Out)
	);
	Batch_Norm bn_kernel26(
		.Data_A(32'b00111110011000000000111001110111),
		.Data_B(32'b00111110101100010001111010111001),
		.Data_In(add_k26_Data_Out),
		.Valid_In(add_kernel26_Valid_Out),
		.Data_Out(bn26_Data_Out),
		.Valid_Out(bn26_Valid_Out)
	);
	Relu_Core rl_kernel26(
		.Data_In(bn26_Data_Out),
		.Valid_In(bn26_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(rl26_Valid_Out)
	);
//////////KERNEL27//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110100001001110110100101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111110000110001011101011001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110111001110111010110001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110100111001111110111100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111101101010011000101101100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110000110101001101101101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111101100111110111111101101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111110110010110011111010100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111110111101110000001101111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111101011111101100001101110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110110111111000110110110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111110100000001011001001000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111111000011011011111100010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111101100001010010001110101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111111011111011010000100101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111110010011110101101100111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111111000011010100000011100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111110111010101010000111010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111110000010000111110011011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110110000100110100000011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111111010110011101001101111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111110101000111101100101111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111110101111001001000110100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111011001101001100010101101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111110100101010111100111010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111110101101101101110110111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111110000011010011110101010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111110010001000000000000111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111111001001010101110000010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111110010101110010110111110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111110001001110011111011111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111100000101111011000001110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel27_Valid_Out)
	);
	Adder_32input add_k27(
		.Data1(Data_Out_Kernel27[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel27[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel27[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel27[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel27[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel27[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel27[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel27[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel27[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel27[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel27[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel27[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel27[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel27[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel27[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel27[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel27[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel27[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel27[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel27[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel27[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel27[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel27[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel27[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel27[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel27[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel27[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel27[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel27[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel27[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel27[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel27[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel27),
		.Data_Out(add_k27_Data_Out),
		.Valid_Out(add_kernel27_Valid_Out)
	);
	Batch_Norm bn_kernel27(
		.Data_A(32'b00111110010101011101001101011110),
		.Data_B(32'b10111110001010101111010100010110),
		.Data_In(add_k27_Data_Out),
		.Valid_In(add_kernel27_Valid_Out),
		.Data_Out(bn27_Data_Out),
		.Valid_Out(bn27_Valid_Out)
	);
	Relu_Core rl_kernel27(
		.Data_In(bn27_Data_Out),
		.Valid_In(bn27_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(rl27_Valid_Out)
	);
//////////KERNEL28//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111101111000110110010000110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111101000110110100111111110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111101101010110100011000111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110100011010101010010101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111101011010100011000000100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111110011110000000010011010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111110101011100101101010001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111110101000100011011000001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111101110110011110011111110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110110001011000100110100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110000110011110001001001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110000111010110100100001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110010111000001110010001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111110001111001000010010101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111101100001111101001111000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111110101001111110101100110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111101111011110000111100010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111110000011100001101110000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111111000011101001001000111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111110110010101110000010010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110101000010100110010010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111111100010000101001110111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110011100111000110110000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111111000111101011011001011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111110100001010000010100101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110000000110111000000001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111110101100000110101001001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111110101100011010100011100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111110111110000011000001101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111111000011110011000111110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111111001101010111010000110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110100100010000110111010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel28_Valid_Out)
	);
	Adder_32input add_k28(
		.Data1(Data_Out_Kernel28[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel28[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel28[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel28[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel28[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel28[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel28[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel28[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel28[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel28[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel28[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel28[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel28[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel28[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel28[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel28[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel28[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel28[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel28[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel28[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel28[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel28[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel28[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel28[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel28[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel28[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel28[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel28[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel28[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel28[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel28[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel28[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel28),
		.Data_Out(add_k28_Data_Out),
		.Valid_Out(add_kernel28_Valid_Out)
	);
	Batch_Norm bn_kernel28(
		.Data_A(32'b00111110010110111000010001000010),
		.Data_B(32'b00111110000010100010011000010100),
		.Data_In(add_k28_Data_Out),
		.Valid_In(add_kernel28_Valid_Out),
		.Data_Out(bn28_Data_Out),
		.Valid_Out(bn28_Valid_Out)
	);
	Relu_Core rl_kernel28(
		.Data_In(bn28_Data_Out),
		.Valid_In(bn28_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(rl28_Valid_Out)
	);
//////////KERNEL29//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111111000110110010101111000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111111100000001110111100111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111111000100001011010110100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110000011110001011010111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111101011101001001011101011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110101101000111110110010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111110100010101100101001000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111110111000110000110001000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111101110011101011000100111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110100101011111110100111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111110000001010011011100101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111100001001100111100110101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111110001000111010011100111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111110001011100000101001111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110111111010001010011110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111110110111011001100100110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111110101001001010001011111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111111011010010000110000010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110100000111010100001111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111101111001001000111111100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110110001000110110111110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111110001000100000111010000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111110001101000110000111111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111110011000001011101101010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111110101100101100100101001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111110100010110111100100110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111110100110110000101110100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111101100000011100110101000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111110110101001011001010000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111101001000000111001010000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111101111000000000100110001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110100001101100111110101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel29_Valid_Out)
	);
	Adder_32input add_k29(
		.Data1(Data_Out_Kernel29[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel29[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel29[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel29[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel29[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel29[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel29[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel29[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel29[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel29[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel29[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel29[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel29[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel29[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel29[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel29[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel29[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel29[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel29[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel29[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel29[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel29[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel29[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel29[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel29[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel29[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel29[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel29[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel29[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel29[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel29[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel29[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel29),
		.Data_Out(add_k29_Data_Out),
		.Valid_Out(add_kernel29_Valid_Out)
	);
	Batch_Norm bn_kernel29(
		.Data_A(32'b00111110100011110001111001111000),
		.Data_B(32'b00111111101000011010100010001111),
		.Data_In(add_k29_Data_Out),
		.Valid_In(add_kernel29_Valid_Out),
		.Data_Out(bn29_Data_Out),
		.Valid_Out(bn29_Valid_Out)
	);
	Relu_Core rl_kernel29(
		.Data_In(bn29_Data_Out),
		.Valid_In(bn29_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(rl29_Valid_Out)
	);
//////////KERNEL30//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111101011011001010100110101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111101011101111111010011001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110010000011001011111110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110010101101000011100110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111111001000110110000001011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111111001011010000010010011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111101011111111110100110100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111101111010000101011111010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111100101010001011001111011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110010101010001011111100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111110101000101111101011001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110101101011000110001100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111111000010000001001101010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111110110001001000001000100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111100100110010010110010110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111110001010000111101001100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111110101101000000100100100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111101100101111111101010101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111110101000100000100011101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110111100111010101011101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110111110101100101110110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111111000110011100001110011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111110100101010011000001011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111111000010011000010100000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111101110100101010100001101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111111000100001101000110100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110001011000100001100000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110000000111110111100100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111111001010000101011110001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110010101100110101000111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111101110000100101100110101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111111001100011110001001111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel30_Valid_Out)
	);
	Adder_32input add_k30(
		.Data1(Data_Out_Kernel30[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel30[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel30[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel30[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel30[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel30[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel30[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel30[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel30[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel30[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel30[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel30[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel30[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel30[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel30[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel30[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel30[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel30[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel30[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel30[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel30[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel30[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel30[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel30[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel30[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel30[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel30[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel30[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel30[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel30[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel30[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel30[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel30),
		.Data_Out(add_k30_Data_Out),
		.Valid_Out(add_kernel30_Valid_Out)
	);
	Batch_Norm bn_kernel30(
		.Data_A(32'b00111110010101110000101011000110),
		.Data_B(32'b00111111001011111110011000110011),
		.Data_In(add_k30_Data_Out),
		.Valid_In(add_kernel30_Valid_Out),
		.Data_Out(bn30_Data_Out),
		.Valid_Out(bn30_Valid_Out)
	);
	Relu_Core rl_kernel30(
		.Data_In(bn30_Data_Out),
		.Valid_In(bn30_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(rl30_Valid_Out)
	);
//////////KERNEL31//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111101110010001111110111010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110101001011011001011000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111101000000100011010001000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111101100001001101110011110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111110110000010001110011100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111100101000101010100101010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111101101000011000011110101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111101000111001001111010110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111100111110101101110000000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110111010110010011001110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111110101101110100011100110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111111000111100100011010010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111110010000100101000010011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111110110110010011110001011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111101110001010010011011110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111110110111011000111010010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111110111010111011111100100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110000110110111100110101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110100111000010111110110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110101001000111001001011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111101100010000010100001110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111110110100000010000100110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110100100111011011100100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111111000011010001100110001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111110010100101101110101100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111111000100100011100010000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111111000101001000100111011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110000100010110100111001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111110001000000111011111101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111111010010110100110110000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111110100100010010001000101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111110111001111101001100001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel31_Valid_Out)
	);
	Adder_32input add_k31(
		.Data1(Data_Out_Kernel31[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel31[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel31[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel31[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel31[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel31[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel31[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel31[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel31[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel31[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel31[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel31[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel31[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel31[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel31[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel31[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel31[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel31[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel31[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel31[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel31[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel31[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel31[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel31[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel31[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel31[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel31[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel31[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel31[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel31[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel31[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel31[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel31),
		.Data_Out(add_k31_Data_Out),
		.Valid_Out(add_kernel31_Valid_Out)
	);
	Batch_Norm bn_kernel31(
		.Data_A(32'b00111110100100010001100100100011),
		.Data_B(32'b00111111110000010011100100011001),
		.Data_In(add_k31_Data_Out),
		.Valid_In(add_kernel31_Valid_Out),
		.Data_Out(bn31_Data_Out),
		.Valid_Out(bn31_Valid_Out)
	);
	Relu_Core rl_kernel31(
		.Data_In(bn31_Data_Out),
		.Valid_In(bn31_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(rl31_Valid_Out)
	);
//////////KERNEL32//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111110101011111000010010001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111100110100110100000001010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110101001001110101110101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110000110010101100111011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111110001000110111011011111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111111000100000100011110100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111110011001100101100110000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111110110111111011000101100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111111100100111111011010001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111111011000110011111100101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110100011010000110000101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111110000100011011000111001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110000001110011011110101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111101110001011011110101111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110010010100000010011000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111110010011101110001110011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111101100110100101001001001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111100101110111111101111011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111110000100001010011111101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111110111000000111100100000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111111001010111111110101000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111101110000001110110110001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111111000110111101000100010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111110011111110110000111000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111110010000001001000010100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111101100001111110001001011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110100010101111011111010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110000111010100101111011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111110101000010011101100100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110001101011100110111011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111101101000011101111010111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110010110010000101010001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel32_Valid_Out)
	);
	Adder_32input add_k32(
		.Data1(Data_Out_Kernel32[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel32[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel32[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel32[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel32[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel32[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel32[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel32[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel32[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel32[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel32[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel32[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel32[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel32[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel32[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel32[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel32[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel32[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel32[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel32[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel32[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel32[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel32[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel32[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel32[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel32[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel32[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel32[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel32[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel32[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel32[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel32[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel32),
		.Data_Out(add_k32_Data_Out),
		.Valid_Out(add_kernel32_Valid_Out)
	);
	Batch_Norm bn_kernel32(
		.Data_A(32'b00111110100111011110011010100100),
		.Data_B(32'b00111101111001010000001011011000),
		.Data_In(add_k32_Data_Out),
		.Valid_In(add_kernel32_Valid_Out),
		.Data_Out(bn32_Data_Out),
		.Valid_Out(bn32_Valid_Out)
	);
	Relu_Core rl_kernel32(
		.Data_In(bn32_Data_Out),
		.Valid_In(bn32_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(rl32_Valid_Out)
	);
//////////KERNEL33//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111110111110110011111011010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111111000001001000110011110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111101101000010011110111000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111101110111100011011011000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111111010111100110000000111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111100010111111111000101100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111110100110101000111000110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111101000001111110000110111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110110100000000110101101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110100001011011100100011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111101110010100010101101000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111101101000001101000000000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111101010000011101011000011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111110000010011000110011000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111111010101110010010010001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111110101000010000001001001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111100101001010101010111110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111101101011000001000110111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111110110010011110010000010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111110110000101101001011111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110000010100100100101001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111111010111010001010111001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110010000010001000010101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111110111100000100101010110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111110101001101100010110101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111111000011011011100110110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110111000001111001101101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110101100010110110101010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111011101011100011111100101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111011000011010000110011010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111110010111111111000010100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111110010001011000001011011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel33_Valid_Out)
	);
	Adder_32input add_k33(
		.Data1(Data_Out_Kernel33[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel33[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel33[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel33[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel33[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel33[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel33[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel33[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel33[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel33[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel33[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel33[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel33[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel33[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel33[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel33[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel33[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel33[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel33[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel33[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel33[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel33[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel33[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel33[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel33[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel33[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel33[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel33[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel33[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel33[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel33[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel33[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel33),
		.Data_Out(add_k33_Data_Out),
		.Valid_Out(add_kernel33_Valid_Out)
	);
	Batch_Norm bn_kernel33(
		.Data_A(32'b00111110010110100100100010000100),
		.Data_B(32'b00111111001101111000010110110000),
		.Data_In(add_k33_Data_Out),
		.Valid_In(add_kernel33_Valid_Out),
		.Data_Out(bn33_Data_Out),
		.Valid_Out(bn33_Valid_Out)
	);
	Relu_Core rl_kernel33(
		.Data_In(bn33_Data_Out),
		.Valid_In(bn33_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(rl33_Valid_Out)
	);
//////////KERNEL34//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111101001011011010100010011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111101100010111100000111101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110100111111011110100110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110111010001011101100010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111110011000010011111111100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111110111101111001010110110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111110101011000101010101100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111101000100010001010001111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111101111101010010011101101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110011010010101011001100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111110000001100010010100011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111110001110001111111001010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110001110000100111011101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111100101011110010111001000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111111010111110011011010101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111110000101010111011100001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111100100111111000000100010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111010101010100110010110111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111111000000010010100101110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111111001100111011111110101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110000000100010100011010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111110111111111100011011010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111111001000101010101011101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111110000100100001000110111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111111001101000001110101100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111100001110000001000001011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110101000011000010001110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110011011111001000001111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111101111100010001100000010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110101000010101110011101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111111000010010010101100110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111101110111111101101001100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel34_Valid_Out)
	);
	Adder_32input add_k34(
		.Data1(Data_Out_Kernel34[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel34[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel34[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel34[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel34[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel34[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel34[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel34[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel34[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel34[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel34[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel34[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel34[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel34[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel34[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel34[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel34[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel34[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel34[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel34[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel34[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel34[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel34[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel34[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel34[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel34[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel34[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel34[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel34[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel34[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel34[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel34[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel34),
		.Data_Out(add_k34_Data_Out),
		.Valid_Out(add_kernel34_Valid_Out)
	);
	Batch_Norm bn_kernel34(
		.Data_A(32'b00111110100000010101001000101000),
		.Data_B(32'b00111111101100110110010101000110),
		.Data_In(add_k34_Data_Out),
		.Valid_In(add_kernel34_Valid_Out),
		.Data_Out(bn34_Data_Out),
		.Valid_Out(bn34_Valid_Out)
	);
	Relu_Core rl_kernel34(
		.Data_In(bn34_Data_Out),
		.Valid_In(bn34_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(rl34_Valid_Out)
	);
//////////KERNEL35//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111101110000000000011111110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111100110111110110001001101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110001101010100011001101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110000000011011011001111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111111000011110000110001000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110010011100011000110111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111111000111101101110000110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111110101101000000011111101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111111100110100010100110000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110101111100000011100110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110111100000010001100000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111100111101100001101111111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110101000010101001101011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111100000011001110001011110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110111011010111110010110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111111000001100000011100100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111110100111010000011110000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110010011100011010101010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111101001010001100011110010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110101101010011011011000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111101000101111000100100001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111110001100001010110010000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110100011010111001111010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111110100110110010011001110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111110111010110011111101101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111110001001011101100111101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110110010010101100100001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110101101001100110010101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111110001110111101110100011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110000111101000001010000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111110110001010100100011111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111110000001001011001000011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel35_Valid_Out)
	);
	Adder_32input add_k35(
		.Data1(Data_Out_Kernel35[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel35[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel35[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel35[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel35[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel35[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel35[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel35[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel35[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel35[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel35[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel35[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel35[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel35[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel35[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel35[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel35[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel35[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel35[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel35[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel35[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel35[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel35[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel35[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel35[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel35[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel35[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel35[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel35[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel35[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel35[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel35[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel35),
		.Data_Out(add_k35_Data_Out),
		.Valid_Out(add_kernel35_Valid_Out)
	);
	Batch_Norm bn_kernel35(
		.Data_A(32'b00111110100101111110110110100111),
		.Data_B(32'b00111111010000010110100110011110),
		.Data_In(add_k35_Data_Out),
		.Valid_In(add_kernel35_Valid_Out),
		.Data_Out(bn35_Data_Out),
		.Valid_Out(bn35_Valid_Out)
	);
	Relu_Core rl_kernel35(
		.Data_In(bn35_Data_Out),
		.Valid_In(bn35_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(rl35_Valid_Out)
	);
//////////KERNEL36//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110100001111011100001100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110101001100100101111001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110100010010000000001110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110001111000100111110011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111111010000010001100110010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110110011100100000011011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111101101010001010000110010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111101100101101010010000000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111110100101011111001000111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111101010101011110110001011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111101010001110000100101001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111110000011101100110111111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110101101100111000001011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111110011010100001010101010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110011001010011101010110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111111000110011110110001011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111101001010000100000010110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111111001101010110100000100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111111100000101110001100110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110110011101111100100111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111111000010110000110011000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111101001000010011000100111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110101010110110001100010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111101110111010011010000010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111101110101000110010010110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111111000011001111010001111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110100001001001011100001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110110111010111101100101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111110100100110010011111101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111011110111001001100010101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111101100011011001010000000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111110001100000110111011010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel36_Valid_Out)
	);
	Adder_32input add_k36(
		.Data1(Data_Out_Kernel36[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel36[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel36[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel36[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel36[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel36[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel36[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel36[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel36[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel36[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel36[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel36[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel36[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel36[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel36[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel36[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel36[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel36[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel36[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel36[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel36[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel36[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel36[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel36[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel36[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel36[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel36[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel36[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel36[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel36[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel36[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel36[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel36),
		.Data_Out(add_k36_Data_Out),
		.Valid_Out(add_kernel36_Valid_Out)
	);
	Batch_Norm bn_kernel36(
		.Data_A(32'b00111110100100100001000000010111),
		.Data_B(32'b00111110011000000111010000111101),
		.Data_In(add_k36_Data_Out),
		.Valid_In(add_kernel36_Valid_Out),
		.Data_Out(bn36_Data_Out),
		.Valid_Out(bn36_Valid_Out)
	);
	Relu_Core rl_kernel36(
		.Data_In(bn36_Data_Out),
		.Valid_In(bn36_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(rl36_Valid_Out)
	);
//////////KERNEL37//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110100011011100011010110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111101101000001101010001011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110101111011011101000110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111111000101101010001011101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111110101001000111000010101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110100010011011101111000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111110001101001110001110000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111101010011110010101110011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111111001011000010001011011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111110100110100000101001011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111100010111000110111011100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111101110110111000110100010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111110100111010010101011011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111101111001001111000001111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110000110001100001011000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111110100011111011111001111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111110011110111010011100110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111101000011101000100100100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110101000110111010100010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110000011111110000000010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111111011010000001100110001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111110110010100101101111001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110110011101111001011010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111111000010101011100001011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111110100111100111100010000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111111000000111100110010010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111111000001101001111100110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110010000011110100001111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111100110001111010010101110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110100001000110100111001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111111000100100011101000000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111110100011001100101101110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel37_Valid_Out)
	);
	Adder_32input add_k37(
		.Data1(Data_Out_Kernel37[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel37[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel37[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel37[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel37[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel37[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel37[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel37[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel37[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel37[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel37[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel37[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel37[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel37[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel37[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel37[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel37[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel37[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel37[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel37[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel37[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel37[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel37[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel37[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel37[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel37[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel37[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel37[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel37[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel37[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel37[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel37[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel37),
		.Data_Out(add_k37_Data_Out),
		.Valid_Out(add_kernel37_Valid_Out)
	);
	Batch_Norm bn_kernel37(
		.Data_A(32'b00111110100100100100100010110000),
		.Data_B(32'b00111111011001110101110010010001),
		.Data_In(add_k37_Data_Out),
		.Valid_In(add_kernel37_Valid_Out),
		.Data_Out(bn37_Data_Out),
		.Valid_Out(bn37_Valid_Out)
	);
	Relu_Core rl_kernel37(
		.Data_In(bn37_Data_Out),
		.Valid_In(bn37_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(rl37_Valid_Out)
	);
//////////KERNEL38//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111010001111101100011010000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111110010110110010001111110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111101101110111100001001101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110000001011001000111101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111110110001101110110111001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111100011001101100000001111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111110110010100110001111110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111110001011101111001001000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110101101000100000000111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110000111110001101100010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111101111100000001010001000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110011110100000100110111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111110100000111001000000011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111110100000110100111000110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110111010100010111000111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111110011010010001000010100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110100000011111011001100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110000010000110001101011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110111001010000010010110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111100100110010100111001111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111111000011001110001111101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111111101010011101001000111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111100010111010010001100001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111110011111100110111010010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111101010100100101011110001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111101101011010110110011100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110110101011101010011000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110001001111100010011011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111111001100100010101000011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110001101011000010001111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111110111000001101111011110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111110101110100010010101110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel38_Valid_Out)
	);
	Adder_32input add_k38(
		.Data1(Data_Out_Kernel38[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel38[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel38[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel38[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel38[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel38[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel38[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel38[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel38[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel38[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel38[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel38[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel38[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel38[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel38[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel38[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel38[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel38[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel38[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel38[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel38[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel38[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel38[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel38[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel38[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel38[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel38[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel38[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel38[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel38[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel38[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel38[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel38),
		.Data_Out(add_k38_Data_Out),
		.Valid_Out(add_kernel38_Valid_Out)
	);
	Batch_Norm bn_kernel38(
		.Data_A(32'b00111110010011101101101101100011),
		.Data_B(32'b00111111001100101001100001101110),
		.Data_In(add_k38_Data_Out),
		.Valid_In(add_kernel38_Valid_Out),
		.Data_Out(bn38_Data_Out),
		.Valid_Out(bn38_Valid_Out)
	);
	Relu_Core rl_kernel38(
		.Data_In(bn38_Data_Out),
		.Valid_In(bn38_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(rl38_Valid_Out)
	);
//////////KERNEL39//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111110010011010010100000100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111110101100011000010010001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110001010100101111011100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110000001001001001110111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111110100010011010111101100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111111001001001100011001001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111110100100010101010001110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111101101111110100010110010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111111000110111001011100110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111101010101110110010101110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111110101111001000001110110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111101110011111011111001000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111110100101010110010110101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111100100101001101010001011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110011110100011111101110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111110111111111111111100101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111110001100111011001001001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111101100111011010110101101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111100100000011101010001010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111101001001010010001010111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111101111000010110001111010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111110010101101110100110010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110110110111011000101001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111111100101000101010110101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111110101100100010111010100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110011110001011010111000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111111001110010000110001111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111111011001011100111100011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111110010000010011011101010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110001011000111101001100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111110010111000110010000011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111110100111100010000100011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel39_Valid_Out)
	);
	Adder_32input add_k39(
		.Data1(Data_Out_Kernel39[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel39[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel39[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel39[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel39[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel39[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel39[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel39[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel39[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel39[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel39[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel39[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel39[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel39[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel39[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel39[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel39[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel39[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel39[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel39[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel39[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel39[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel39[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel39[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel39[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel39[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel39[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel39[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel39[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel39[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel39[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel39[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel39),
		.Data_Out(add_k39_Data_Out),
		.Valid_Out(add_kernel39_Valid_Out)
	);
	Batch_Norm bn_kernel39(
		.Data_A(32'b00111110011100011011001010010000),
		.Data_B(32'b00111111001000110110101000000100),
		.Data_In(add_k39_Data_Out),
		.Valid_In(add_kernel39_Valid_Out),
		.Data_Out(bn39_Data_Out),
		.Valid_Out(bn39_Valid_Out)
	);
	Relu_Core rl_kernel39(
		.Data_In(bn39_Data_Out),
		.Valid_In(bn39_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(rl39_Valid_Out)
	);
//////////KERNEL40//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111101100000111011011001001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110000101000111010100010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111100110000001000001000010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110100101100000010111100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111101001111100111011001000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111101000111110101111110100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111110100001010110100010111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111101100001110100101110000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111101101011001110001001101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110011000010001110110101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111111001001100001101001001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111101110111100010100100010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111101111010101111111100100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111110011010101010000100110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111101010001001111000001100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111101001001010000100110100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111111000100110110101011001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111101101111000100100001100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111110100000111000101111101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111111000101111101011001100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111111000100110001010000010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111101011110010001101010010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111111010011100001000011001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111110100100000001111010111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111110100111010100110010000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111111011101101000101000001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111111000011001111001101101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111100101110001011111000000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111110100100010000000110110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111101000001111011110111011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111110100000100101000011000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111111010000000101110101001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel40_Valid_Out)
	);
	Adder_32input add_k40(
		.Data1(Data_Out_Kernel40[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel40[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel40[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel40[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel40[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel40[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel40[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel40[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel40[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel40[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel40[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel40[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel40[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel40[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel40[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel40[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel40[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel40[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel40[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel40[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel40[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel40[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel40[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel40[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel40[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel40[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel40[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel40[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel40[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel40[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel40[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel40[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel40),
		.Data_Out(add_k40_Data_Out),
		.Valid_Out(add_kernel40_Valid_Out)
	);
	Batch_Norm bn_kernel40(
		.Data_A(32'b00111110011111111001001001001100),
		.Data_B(32'b10111111001101101000011011111100),
		.Data_In(add_k40_Data_Out),
		.Valid_In(add_kernel40_Valid_Out),
		.Data_Out(bn40_Data_Out),
		.Valid_Out(bn40_Valid_Out)
	);
	Relu_Core rl_kernel40(
		.Data_In(bn40_Data_Out),
		.Valid_In(bn40_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(rl40_Valid_Out)
	);
//////////KERNEL41//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111111000110111000010001001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111110100111100111101101010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111101010100111101100000110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111101010111101000111111100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111111010010011011100000010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111111001010001001011011111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111110001000101110101111001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111110010000001001010010111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110010011000101010011110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110110101001111111111101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111111010010001110010111110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110011011111110001001000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110111001010001101001001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111110110011011111100010010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111101011101000011100110111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111101101011000111001011110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111110011100000100100010011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111110010010000101101110110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110101101000011010110110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111110111111100111001100000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110110011000010000110001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111011100001010100101100101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110101100101001001100101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111111001101001001100101101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111100111100110011111100110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110110100111000111100110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111110110000101000111111101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111110100010100111000111011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111110000101111100011111011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110001011111111110110001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111100010110110111101111000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111101011101100101110000010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel41_Valid_Out)
	);
	Adder_32input add_k41(
		.Data1(Data_Out_Kernel41[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel41[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel41[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel41[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel41[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel41[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel41[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel41[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel41[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel41[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel41[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel41[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel41[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel41[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel41[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel41[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel41[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel41[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel41[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel41[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel41[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel41[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel41[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel41[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel41[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel41[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel41[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel41[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel41[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel41[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel41[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel41[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel41),
		.Data_Out(add_k41_Data_Out),
		.Valid_Out(add_kernel41_Valid_Out)
	);
	Batch_Norm bn_kernel41(
		.Data_A(32'b00111110101010010001111010101000),
		.Data_B(32'b00111111000101000101110101111111),
		.Data_In(add_k41_Data_Out),
		.Valid_In(add_kernel41_Valid_Out),
		.Data_Out(bn41_Data_Out),
		.Valid_Out(bn41_Valid_Out)
	);
	Relu_Core rl_kernel41(
		.Data_In(bn41_Data_Out),
		.Valid_In(bn41_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(rl41_Valid_Out)
	);
//////////KERNEL42//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111110111010110010110001111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111101011001010101110101010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110001000000000110100110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110011100100011010000000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111111000010010001110000011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110001110100110110000010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111101101001001110011010010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111101000001111010110111011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110000010000000110001011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111110110110111101011100110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111111000000011001111001011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111101101011010111001000000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111101100001000101010000011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111100110011100100100010011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110101000100001100011001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111110010010000001111010110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111110001001110001001001110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111101110101110001000110110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110000110101001100101100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111110000111010111001110001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111111100100000001001011000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111110011001010001000001001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111110100001010100100011110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111010011001111010000010111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111111001000100100010111101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111111001011111110100000011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111110110101011001101010111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110101000010001110010111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111110101110111011110110111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110111110011001101100011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111101100000101011000101100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111110100101000011011000000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel42_Valid_Out)
	);
	Adder_32input add_k42(
		.Data1(Data_Out_Kernel42[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel42[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel42[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel42[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel42[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel42[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel42[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel42[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel42[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel42[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel42[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel42[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel42[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel42[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel42[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel42[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel42[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel42[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel42[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel42[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel42[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel42[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel42[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel42[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel42[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel42[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel42[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel42[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel42[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel42[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel42[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel42[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel42),
		.Data_Out(add_k42_Data_Out),
		.Valid_Out(add_kernel42_Valid_Out)
	);
	Batch_Norm bn_kernel42(
		.Data_A(32'b00111110100010101100100100110101),
		.Data_B(32'b00111111001010110010101001000101),
		.Data_In(add_k42_Data_Out),
		.Valid_In(add_kernel42_Valid_Out),
		.Data_Out(bn42_Data_Out),
		.Valid_Out(bn42_Valid_Out)
	);
	Relu_Core rl_kernel42(
		.Data_In(bn42_Data_Out),
		.Valid_In(bn42_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(rl42_Valid_Out)
	);
//////////KERNEL43//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110101100011011111111110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110100111000100100011000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110111011000101000011001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111101001100000100110000110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111110001001001101100001011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110100111100010100100001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111110001011101110111110101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111101011110010001010000111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111110111110110110110011010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110101111001111111110001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111110110101111010000010101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110111000101011110010000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110001011101100001111010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111110110111001011000010011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110011011111110110010010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111101100111001001110001101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111111000011111001100100000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111101100101011011101101100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110110100100100001010110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110010001110100011111110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110110100011011100111001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111110110000011001101101010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111100110001100001100010101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111111010110010001101101010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111100110100001001101101100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111110111110011110000011100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111110001001001011010001011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111110100001101011101110101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111110110000110001011011101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111101110110000100010001000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111101001111110011100101110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111111001100110011111000001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel43_Valid_Out)
	);
	Adder_32input add_k43(
		.Data1(Data_Out_Kernel43[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel43[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel43[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel43[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel43[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel43[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel43[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel43[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel43[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel43[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel43[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel43[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel43[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel43[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel43[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel43[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel43[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel43[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel43[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel43[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel43[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel43[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel43[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel43[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel43[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel43[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel43[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel43[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel43[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel43[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel43[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel43[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel43),
		.Data_Out(add_k43_Data_Out),
		.Valid_Out(add_kernel43_Valid_Out)
	);
	Batch_Norm bn_kernel43(
		.Data_A(32'b00111110111010100000011101011010),
		.Data_B(32'b00111111011111001000011001010101),
		.Data_In(add_k43_Data_Out),
		.Valid_In(add_kernel43_Valid_Out),
		.Data_Out(bn43_Data_Out),
		.Valid_Out(bn43_Valid_Out)
	);
	Relu_Core rl_kernel43(
		.Data_In(bn43_Data_Out),
		.Valid_In(bn43_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(rl43_Valid_Out)
	);
//////////KERNEL44//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111101011101110001101101100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111111010011010111010001101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110100001100010001001001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110101110000100011111010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111110000010101001000110011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110110010110000100000000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111110100010111100110110101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111011000001110101110101011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110101110011111000110110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111110011100010001111100110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110110110101110000101100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110010101110111010101101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111101101100101100111101011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111111000101000000111101010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110110010011011001110010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111110000001010001001111111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111110100111001100101111111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110111001110001010111001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110101100011100010100000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111101111011111011011001111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110100010101100111011111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111110100110011101000011110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110101001101001111100011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111110100100000110110011000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111111001101111011000000100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111101111110011110000111111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110000000111001010101000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110101010010011001110100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111111000010001101010000011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110101011111000101100110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111110110000000111100100011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110010101111111001000101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel44_Valid_Out)
	);
	Adder_32input add_k44(
		.Data1(Data_Out_Kernel44[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel44[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel44[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel44[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel44[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel44[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel44[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel44[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel44[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel44[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel44[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel44[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel44[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel44[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel44[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel44[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel44[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel44[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel44[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel44[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel44[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel44[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel44[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel44[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel44[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel44[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel44[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel44[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel44[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel44[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel44[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel44[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel44),
		.Data_Out(add_k44_Data_Out),
		.Valid_Out(add_kernel44_Valid_Out)
	);
	Batch_Norm bn_kernel44(
		.Data_A(32'b00111110101000110111001001011100),
		.Data_B(32'b00111111100001100110110111111000),
		.Data_In(add_k44_Data_Out),
		.Valid_In(add_kernel44_Valid_Out),
		.Data_Out(bn44_Data_Out),
		.Valid_Out(bn44_Valid_Out)
	);
	Relu_Core rl_kernel44(
		.Data_In(bn44_Data_Out),
		.Valid_In(bn44_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(rl44_Valid_Out)
	);
//////////KERNEL45//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111111000010011100100101101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111110010011011000011101000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110100001101111110110111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110001110001010110000111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111101110011010001001110010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110000110001111101001101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111101100000100000001000110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111100000011111101110000000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111110111111100000001010110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110001111000011001101000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111110001100110110110001100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111110000110101100100010011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111101111011000110101001111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111101001000100011101110010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110011000011110110000010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111110111010010000001101101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111101111101010101011000011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110101000110100010101100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110000000001001110110101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111111011111110111010111100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111111000100100111000010011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111110101111000110101001011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111101101110010001101011001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111110100111111111010101110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111111001001000001001101001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111100111111110001111001100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111101011100101000010000011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111101100010111111111010101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111110111100000010010000000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111111000011011010100101110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111110111110011100100110111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111111000010100100011000011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel45_Valid_Out)
	);
	Adder_32input add_k45(
		.Data1(Data_Out_Kernel45[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel45[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel45[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel45[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel45[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel45[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel45[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel45[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel45[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel45[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel45[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel45[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel45[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel45[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel45[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel45[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel45[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel45[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel45[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel45[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel45[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel45[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel45[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel45[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel45[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel45[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel45[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel45[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel45[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel45[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel45[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel45[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel45),
		.Data_Out(add_k45_Data_Out),
		.Valid_Out(add_kernel45_Valid_Out)
	);
	Batch_Norm bn_kernel45(
		.Data_A(32'b00111110101010011010001101111101),
		.Data_B(32'b00111110101111011000011011111101),
		.Data_In(add_k45_Data_Out),
		.Valid_In(add_kernel45_Valid_Out),
		.Data_Out(bn45_Data_Out),
		.Valid_Out(bn45_Valid_Out)
	);
	Relu_Core rl_kernel45(
		.Data_In(bn45_Data_Out),
		.Valid_In(bn45_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(rl45_Valid_Out)
	);
//////////KERNEL46//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111111000010000001001010100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111110111001110011000001000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110101110010000010010000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111111010101110111110101101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111110100101000001011110101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110000100110101010001101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111110010000011000001010011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111110011101101100110010010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111111000001100111111011010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111101110100000101101000011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110111000100010010011011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111111001111101100101101111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111101100101101110011110000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111110010110100011101001000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110100001111101011110111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111110011001000010110110101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111111000001000010010101001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111101000101110001101101011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110010110100110100001011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111110100000011010100111010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110010010000111111111111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111110100101100000001101011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111110000001110110111101110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111110110110000110011100111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111101010111101010011101010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111101010100011010101100000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110011100010110000111001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110100110111100000001000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111101101000001000100110110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111110010010100010000001010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111110111100001101001011011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111101111011001111000000010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel46_Valid_Out)
	);
	Adder_32input add_k46(
		.Data1(Data_Out_Kernel46[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel46[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel46[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel46[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel46[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel46[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel46[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel46[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel46[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel46[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel46[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel46[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel46[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel46[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel46[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel46[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel46[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel46[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel46[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel46[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel46[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel46[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel46[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel46[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel46[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel46[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel46[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel46[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel46[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel46[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel46[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel46[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel46),
		.Data_Out(add_k46_Data_Out),
		.Valid_Out(add_kernel46_Valid_Out)
	);
	Batch_Norm bn_kernel46(
		.Data_A(32'b00111110100001111100101000100011),
		.Data_B(32'b00111110001000010101111010010110),
		.Data_In(add_k46_Data_Out),
		.Valid_In(add_kernel46_Valid_Out),
		.Data_Out(bn46_Data_Out),
		.Valid_Out(bn46_Valid_Out)
	);
	Relu_Core rl_kernel46(
		.Data_In(bn46_Data_Out),
		.Valid_In(bn46_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(rl46_Valid_Out)
	);
//////////KERNEL47//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111111001111000110000010110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111110010100011001100001010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111111001011011000010110110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110110000001100010000001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111101010100101010111000100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111101111001101011100000101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111101001111101010010101000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111110100010000010001100101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111101000101000011101011010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110111010110010110111110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110101101010001111100110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111100111001010110011000100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110110001001110010000110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111011111111010101001000001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110011011000010110110001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111101101010010010010111100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111110011110110010101110101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111110100011011110101001110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111001110111100001011001111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111111000011111111111111011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111111000000101100001110011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111110011001001101000100011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110101010100010000001110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111111000000001100000001110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111111010010101100100000100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111111000110000010010111001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111110101010101011101011001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111100101000011110100111101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111110100001110001010000100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111110000001101001000110011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111111001010000001001000010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110100011000111111101100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel47_Valid_Out)
	);
	Adder_32input add_k47(
		.Data1(Data_Out_Kernel47[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel47[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel47[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel47[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel47[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel47[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel47[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel47[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel47[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel47[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel47[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel47[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel47[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel47[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel47[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel47[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel47[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel47[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel47[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel47[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel47[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel47[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel47[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel47[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel47[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel47[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel47[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel47[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel47[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel47[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel47[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel47[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel47),
		.Data_Out(add_k47_Data_Out),
		.Valid_Out(add_kernel47_Valid_Out)
	);
	Batch_Norm bn_kernel47(
		.Data_A(32'b00111110010010000000110111001010),
		.Data_B(32'b10111110110010000111100111000111),
		.Data_In(add_k47_Data_Out),
		.Valid_In(add_kernel47_Valid_Out),
		.Data_Out(bn47_Data_Out),
		.Valid_Out(bn47_Valid_Out)
	);
	Relu_Core rl_kernel47(
		.Data_In(bn47_Data_Out),
		.Valid_In(bn47_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(rl47_Valid_Out)
	);
//////////KERNEL48//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110000011110110110100110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110110000100110001001111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110000011101011000110101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110101011001011100101001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111110001011001010010110110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111111000111101011001111000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111101111001001101100111111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111110101010001111100001000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111101101110010001000011000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110001010100111110011101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111100110001100000110000000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111110001000100100001110111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110100111111110111000000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111101000000100000110110000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110101101011010011010110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111101111111110111111110111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111110010001000010110110010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111110011111001010010100101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110111100101101000010000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111110101101110101101111011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110101001001110100001110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111111000110100001010001011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110100001010101001101111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111101111011110110001001011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111111000000101010110110101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111110011000110111110100001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111110010010001000010100110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111101101101110011001000000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111111000101101000101110100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111111000000110101100001110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111111010001011010110010111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111111000100000111010000110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel48_Valid_Out)
	);
	Adder_32input add_k48(
		.Data1(Data_Out_Kernel48[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel48[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel48[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel48[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel48[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel48[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel48[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel48[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel48[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel48[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel48[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel48[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel48[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel48[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel48[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel48[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel48[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel48[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel48[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel48[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel48[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel48[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel48[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel48[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel48[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel48[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel48[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel48[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel48[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel48[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel48[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel48[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel48),
		.Data_Out(add_k48_Data_Out),
		.Valid_Out(add_kernel48_Valid_Out)
	);
	Batch_Norm bn_kernel48(
		.Data_A(32'b00111110010111101001011001111100),
		.Data_B(32'b00111110100000101011101110010001),
		.Data_In(add_k48_Data_Out),
		.Valid_In(add_kernel48_Valid_Out),
		.Data_Out(bn48_Data_Out),
		.Valid_Out(bn48_Valid_Out)
	);
	Relu_Core rl_kernel48(
		.Data_In(bn48_Data_Out),
		.Valid_In(bn48_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(rl48_Valid_Out)
	);
//////////KERNEL49//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111111000101100100111010011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111110011001101111010001111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111100111011111010100100110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111101101000111111010000000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111101111000110000011111111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110000000100010001101111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111110110100111110000010001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111110101011000000101111100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111111011100001010100011101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111011010011010001001110001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110111110011110001011010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110000100000011111101111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110011001110001101101000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111101100110000011001010010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111111100111011000111010010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111110001111000011011111010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111110100101100100000001100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111110010011111010010101100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110111011100010110110000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111101001000000111101100101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110001001101011110111110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111110010111110000101010110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111110110000010100000010010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111110000010000111100000010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111110111001001111001100101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111101100010000000110010011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110011110110110111100001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110011011000001101101001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111110100010011111100000011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111110000010100110110101110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111110111000000110011110000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111100010001111110100001111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel49_Valid_Out)
	);
	Adder_32input add_k49(
		.Data1(Data_Out_Kernel49[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel49[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel49[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel49[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel49[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel49[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel49[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel49[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel49[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel49[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel49[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel49[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel49[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel49[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel49[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel49[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel49[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel49[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel49[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel49[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel49[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel49[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel49[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel49[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel49[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel49[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel49[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel49[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel49[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel49[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel49[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel49[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel49),
		.Data_Out(add_k49_Data_Out),
		.Valid_Out(add_kernel49_Valid_Out)
	);
	Batch_Norm bn_kernel49(
		.Data_A(32'b00111110101001001010011100000011),
		.Data_B(32'b10111110000010010100100010110001),
		.Data_In(add_k49_Data_Out),
		.Valid_In(add_kernel49_Valid_Out),
		.Data_Out(bn49_Data_Out),
		.Valid_Out(bn49_Valid_Out)
	);
	Relu_Core rl_kernel49(
		.Data_In(bn49_Data_Out),
		.Valid_In(bn49_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(rl49_Valid_Out)
	);
//////////KERNEL50//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110000110011011010111100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111101010011111010110100000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111111001111101110000110110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110001100001001100000000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111110000001101100001100011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111110111011111110100000101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111110000001010001100100110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111110100001000100111000100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111111001100110011100111000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110110101110011010110111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110111100101010110001111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110011101110010111101100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111101100000011111110010011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111100000111001001110011110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110001000110001011010011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111100111010001000010111010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111110010010001010100100011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110101111111111011001001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111110000110110011011000101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111111000010011100011000000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110000101001001001100001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111001011000001000011110010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111110000100101001100000011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111111000100111010100010111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111110000000111100101100101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110111001110110110110100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110101100110110010010101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111110010011011000101111000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111110111110010110111011000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111110000110000100100110101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111111011110101100111111111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110001100111001001110110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel50_Valid_Out)
	);
	Adder_32input add_k50(
		.Data1(Data_Out_Kernel50[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel50[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel50[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel50[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel50[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel50[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel50[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel50[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel50[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel50[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel50[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel50[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel50[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel50[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel50[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel50[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel50[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel50[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel50[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel50[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel50[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel50[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel50[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel50[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel50[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel50[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel50[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel50[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel50[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel50[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel50[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel50[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel50),
		.Data_Out(add_k50_Data_Out),
		.Valid_Out(add_kernel50_Valid_Out)
	);
	Batch_Norm bn_kernel50(
		.Data_A(32'b00111110011111001000011110001111),
		.Data_B(32'b00111111011001000010000100001111),
		.Data_In(add_k50_Data_Out),
		.Valid_In(add_kernel50_Valid_Out),
		.Data_Out(bn50_Data_Out),
		.Valid_Out(bn50_Valid_Out)
	);
	Relu_Core rl_kernel50(
		.Data_In(bn50_Data_Out),
		.Valid_In(bn50_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(rl50_Valid_Out)
	);
//////////KERNEL51//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111111001000101001011111000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110010111100000110111001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110000001101111110010011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110011110100101100001100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111111011000101000000011000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111101100000011101010010011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111100011000111000111100110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111111000000010001111000111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111101011100001011110110010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110101101001111101011100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111101100001001110000101010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111100101010100011111111100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110001000011111100001000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111111001001101111000001010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110101011010110011000101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111110011001001011001001100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111110001001100111100111100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111110001011001011100110110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111111000100011000000010111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111110000101001100100011010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111101101000001111010010100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111101100010010011111110010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111100101010011011101100100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111110011011000010000100010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111101110010011110101101001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110111101111000011010000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110010110001001010100001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111111100000011010001010100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111101101001100000110111110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111111000011110111111001101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111101101110010110011000010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111110100111001110001101110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel51_Valid_Out)
	);
	Adder_32input add_k51(
		.Data1(Data_Out_Kernel51[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel51[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel51[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel51[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel51[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel51[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel51[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel51[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel51[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel51[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel51[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel51[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel51[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel51[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel51[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel51[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel51[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel51[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel51[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel51[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel51[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel51[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel51[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel51[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel51[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel51[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel51[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel51[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel51[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel51[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel51[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel51[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel51),
		.Data_Out(add_k51_Data_Out),
		.Valid_Out(add_kernel51_Valid_Out)
	);
	Batch_Norm bn_kernel51(
		.Data_A(32'b00111110101100001000100011011001),
		.Data_B(32'b00111111101000010100111100111011),
		.Data_In(add_k51_Data_Out),
		.Valid_In(add_kernel51_Valid_Out),
		.Data_Out(bn51_Data_Out),
		.Valid_Out(bn51_Valid_Out)
	);
	Relu_Core rl_kernel51(
		.Data_In(bn51_Data_Out),
		.Valid_In(bn51_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(rl51_Valid_Out)
	);
//////////KERNEL52//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111111000001000101010100111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111111000000100110001010111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110010110011101110000101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110001001111000001111000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111101010100001011110011011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110001000110010010110001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111110101000111001100100011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111110000101010000100111010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111111011011111101101010011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110100000011111000011000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110100000100011011111111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111101100111001000001110110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110101110111011011101110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111110010100001101110111000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110111111001000110000101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111111000001000010001111001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111110011111111110101001111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111110100010011100011101100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111100100111000001010011100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111101001000000100111010010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110100011101000010001100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111110001111010100110010100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110010111101101111100100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111110100100101100011001110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111101000111010110110010111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111111010110101101011011000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111101001110110110000000001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111110110000001111001000100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111101100010000011000100010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111110000011001011110100100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111110111101101010110011011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111111010001011001110110111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel52_Valid_Out)
	);
	Adder_32input add_k52(
		.Data1(Data_Out_Kernel52[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel52[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel52[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel52[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel52[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel52[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel52[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel52[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel52[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel52[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel52[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel52[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel52[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel52[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel52[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel52[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel52[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel52[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel52[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel52[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel52[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel52[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel52[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel52[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel52[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel52[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel52[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel52[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel52[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel52[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel52[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel52[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel52),
		.Data_Out(add_k52_Data_Out),
		.Valid_Out(add_kernel52_Valid_Out)
	);
	Batch_Norm bn_kernel52(
		.Data_A(32'b00111110011000000111010001001101),
		.Data_B(32'b10111110010010111111011111110001),
		.Data_In(add_k52_Data_Out),
		.Valid_In(add_kernel52_Valid_Out),
		.Data_Out(bn52_Data_Out),
		.Valid_Out(bn52_Valid_Out)
	);
	Relu_Core rl_kernel52(
		.Data_In(bn52_Data_Out),
		.Valid_In(bn52_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(rl52_Valid_Out)
	);
//////////KERNEL53//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111110010000001011111100010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111110001010000010100111100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110110100111111111010000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111101010111100101100000010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111110110011111000011010101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111110001000110000001010011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111101110011000100111100011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111110000110101110110110000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110110110100100010101111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110010000100001011110011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111101011010010110001000110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111101100010000001100000010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110101100011010110011010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111101101111000000010010111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110101111011000110110000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111110110000000111111111101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110101010000011001000101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111110100101001000010011110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110011111011011010111110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111110111011110101000111100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110111010011011010101100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111101011101100011110001000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111110000010101011001010010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111110101010111010110000111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111101110000101001000111011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110111101001000110000111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111111100000011010011110010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110101010001101100101111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111110011110001111000100001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111111000010100000010010010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111101100000011010000001011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111111100000011001100010010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel53_Valid_Out)
	);
	Adder_32input add_k53(
		.Data1(Data_Out_Kernel53[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel53[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel53[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel53[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel53[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel53[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel53[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel53[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel53[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel53[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel53[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel53[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel53[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel53[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel53[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel53[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel53[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel53[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel53[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel53[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel53[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel53[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel53[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel53[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel53[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel53[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel53[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel53[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel53[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel53[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel53[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel53[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel53),
		.Data_Out(add_k53_Data_Out),
		.Valid_Out(add_kernel53_Valid_Out)
	);
	Batch_Norm bn_kernel53(
		.Data_A(32'b00111110100011100100111110100000),
		.Data_B(32'b00111111010110001100100011101111),
		.Data_In(add_k53_Data_Out),
		.Valid_In(add_kernel53_Valid_Out),
		.Data_Out(bn53_Data_Out),
		.Valid_Out(bn53_Valid_Out)
	);
	Relu_Core rl_kernel53(
		.Data_In(bn53_Data_Out),
		.Valid_In(bn53_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(rl53_Valid_Out)
	);
//////////KERNEL54//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110111001001010001101110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110010100000111100010011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111111010111101100001000110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110011000010110101011100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111110110001011101001001111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111110101001110110001011011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111110010001100100111110010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111111000010101111100001001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111111000100000010010111101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111100011011001010100000010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110011010000110110001010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110000111000000111000110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110000100010100100011011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111110000110100001000011010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110101011100100100001111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111111001010011100111110011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111101101001100101001011101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111110111011100101011001100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111101011001000010000010110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111110100111001001111011001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110110110011100010000111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111100111001101100001110010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111110100000000100111011100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111110000101111111111010100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111100001100110000001110111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111101111010100010111110111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110100000111001101101100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111111000110010011100011011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111110101000011001001001110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110111100010011111110101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111110111101110110100111101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110101111000111000001100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel54_Valid_Out)
	);
	Adder_32input add_k54(
		.Data1(Data_Out_Kernel54[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel54[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel54[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel54[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel54[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel54[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel54[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel54[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel54[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel54[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel54[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel54[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel54[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel54[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel54[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel54[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel54[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel54[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel54[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel54[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel54[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel54[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel54[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel54[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel54[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel54[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel54[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel54[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel54[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel54[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel54[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel54[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel54),
		.Data_Out(add_k54_Data_Out),
		.Valid_Out(add_kernel54_Valid_Out)
	);
	Batch_Norm bn_kernel54(
		.Data_A(32'b00111110011001111011001001001000),
		.Data_B(32'b00111111011011110100011111100100),
		.Data_In(add_k54_Data_Out),
		.Valid_In(add_kernel54_Valid_Out),
		.Data_Out(bn54_Data_Out),
		.Valid_Out(bn54_Valid_Out)
	);
	Relu_Core rl_kernel54(
		.Data_In(bn54_Data_Out),
		.Valid_In(bn54_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(rl54_Valid_Out)
	);
//////////KERNEL55//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110001110100111111001010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110100111100111111101101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110101001000001111000110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110101100000000100000100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111110011000100111100000000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111110000010101110101001000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111101001010000010101001001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111110100001111010101111111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110010101110010101111011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110110000101011001000111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110110100010111111100111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110000000000001100000010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111111011010000100011001100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111110101010001011010010101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110110011000000111100011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111110101010110011010111100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111111000101101100110010010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110111000100000000110110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110100001010010000001011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111101101101110111001001000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110111101001011110111011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111101100110100001010011111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111101100100010111001011001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111110111001111000001101011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111111000000100000111111001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111101100011000100010000011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110001100011000010010111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111111000011010110110001010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111110110111000010101010001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110001110101111001000111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111110110001011111001001111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110111001111111100111000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel55_Valid_Out)
	);
	Adder_32input add_k55(
		.Data1(Data_Out_Kernel55[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel55[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel55[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel55[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel55[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel55[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel55[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel55[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel55[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel55[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel55[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel55[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel55[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel55[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel55[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel55[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel55[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel55[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel55[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel55[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel55[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel55[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel55[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel55[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel55[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel55[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel55[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel55[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel55[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel55[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel55[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel55[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel55),
		.Data_Out(add_k55_Data_Out),
		.Valid_Out(add_kernel55_Valid_Out)
	);
	Batch_Norm bn_kernel55(
		.Data_A(32'b00111110011001101101111011000001),
		.Data_B(32'b00111111010000100001011110110101),
		.Data_In(add_k55_Data_Out),
		.Valid_In(add_kernel55_Valid_Out),
		.Data_Out(bn55_Data_Out),
		.Valid_Out(bn55_Valid_Out)
	);
	Relu_Core rl_kernel55(
		.Data_In(bn55_Data_Out),
		.Valid_In(bn55_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(rl55_Valid_Out)
	);
//////////KERNEL56//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111111010101001010011110100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111100111010010100000100000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111101101111101010001000001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110101001101101101001111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111110110100111001000100111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110001001000110001111110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111110101000011110011010100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111110111100000011011101011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110001100010110100010111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111110010100011011000110100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111111000000101101110010001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111110110010010101101011111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110101111111111101110110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111110010101101101000000100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111101111000101000111001110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111111000011101101100100101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111110110111100101111100110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111100101101101101010011000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110011011111001010110010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111111010001011001100100110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111101110000011000001011101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111110101101110011100101100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111110101011100111110111001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111101111000101010000000010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111101111010011010110101000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110110111100000001110010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111110000011110101010000010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111101000010111100101010010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111110011010011010100111010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111101000000011111011101100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111111001010111011111011110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110001011110110110100001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel56_Valid_Out)
	);
	Adder_32input add_k56(
		.Data1(Data_Out_Kernel56[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel56[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel56[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel56[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel56[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel56[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel56[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel56[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel56[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel56[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel56[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel56[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel56[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel56[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel56[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel56[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel56[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel56[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel56[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel56[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel56[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel56[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel56[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel56[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel56[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel56[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel56[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel56[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel56[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel56[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel56[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel56[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel56),
		.Data_Out(add_k56_Data_Out),
		.Valid_Out(add_kernel56_Valid_Out)
	);
	Batch_Norm bn_kernel56(
		.Data_A(32'b00111110100001100111010101110110),
		.Data_B(32'b00111111001011111011000010101100),
		.Data_In(add_k56_Data_Out),
		.Valid_In(add_kernel56_Valid_Out),
		.Data_Out(bn56_Data_Out),
		.Valid_Out(bn56_Valid_Out)
	);
	Relu_Core rl_kernel56(
		.Data_In(bn56_Data_Out),
		.Valid_In(bn56_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(rl56_Valid_Out)
	);
//////////KERNEL57//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110110011100111001000010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110011000011111100111000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110100100011001110001001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110011100000011110011011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111110010010111011010011110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110100011111101111000110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111110000111001001001001010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111110101110101011011000111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111110110000111101110001010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111101101001100111001101010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111110100001110010011000101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110100111011001001000111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110110010111010000110100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111110000101110101110000011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111111001101000010001000000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111110010000011100111001010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111100011111011010101100011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111110000100001000010100000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110010110101111011101000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110111111111011000000111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111101111101000111111001110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111111001010001000101000000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111101111011111100110100111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111110101010011100011111000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111110000000101101010110111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110011111101010001010011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111111100000010000111000001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110100001101101001010010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111110101010111001100011110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110101010011101001010101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111110100011000110001010011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111111001010111100001010111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel57_Valid_Out)
	);
	Adder_32input add_k57(
		.Data1(Data_Out_Kernel57[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel57[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel57[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel57[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel57[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel57[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel57[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel57[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel57[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel57[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel57[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel57[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel57[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel57[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel57[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel57[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel57[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel57[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel57[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel57[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel57[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel57[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel57[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel57[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel57[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel57[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel57[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel57[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel57[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel57[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel57[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel57[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel57),
		.Data_Out(add_k57_Data_Out),
		.Valid_Out(add_kernel57_Valid_Out)
	);
	Batch_Norm bn_kernel57(
		.Data_A(32'b00111110100000101100110110001011),
		.Data_B(32'b00111111011011101010101101011100),
		.Data_In(add_k57_Data_Out),
		.Valid_In(add_kernel57_Valid_Out),
		.Data_Out(bn57_Data_Out),
		.Valid_Out(bn57_Valid_Out)
	);
	Relu_Core rl_kernel57(
		.Data_In(bn57_Data_Out),
		.Valid_In(bn57_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(rl57_Valid_Out)
	);
//////////KERNEL58//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111111011101010110000111110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111011100000100101101101111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111111000001000000111100001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111101110010111011101101101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111101000001111111111100000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110110100111110111000011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111110011111100001001111010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111110101001010111111011001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111101111001110000100110111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110100110011101101001001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111110100001110110011100001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111111000000011010100000011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110101001110011100101111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111110001001010001010001110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110010111001110001111000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111110111101101110100110100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111111001100111101011000000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111110010010010010110110000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110100101100111110001010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111110000110000110001110100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111101100000101101110101010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111110110111010001100001010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110100011001100101011100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111101010100000001011110101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111110101111100001011000000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111101110111111111101111001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110000010001010000000101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111111000000011011000011010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111110110110111011101010011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110110001111000101011011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111100100001000011010101010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111111001000011101010110111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel58_Valid_Out)
	);
	Adder_32input add_k58(
		.Data1(Data_Out_Kernel58[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel58[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel58[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel58[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel58[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel58[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel58[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel58[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel58[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel58[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel58[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel58[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel58[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel58[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel58[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel58[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel58[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel58[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel58[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel58[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel58[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel58[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel58[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel58[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel58[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel58[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel58[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel58[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel58[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel58[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel58[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel58[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel58),
		.Data_Out(add_k58_Data_Out),
		.Valid_Out(add_kernel58_Valid_Out)
	);
	Batch_Norm bn_kernel58(
		.Data_A(32'b00111110010010011001100001101010),
		.Data_B(32'b00111111000011111111000100101011),
		.Data_In(add_k58_Data_Out),
		.Valid_In(add_kernel58_Valid_Out),
		.Data_Out(bn58_Data_Out),
		.Valid_Out(bn58_Valid_Out)
	);
	Relu_Core rl_kernel58(
		.Data_In(bn58_Data_Out),
		.Valid_In(bn58_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(rl58_Valid_Out)
	);
//////////KERNEL59//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111110110110111001011111001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110100110001100101000110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110000011100111000111000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110100000010001001110001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111101010110011100110101000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111101010010000000001000100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111100110001011011100110101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111111001011111111011100111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111101100000101011000100111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111110110011110011000000000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111111001110000000100111001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111101011001001101010001110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111111100001101010000000011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111111000010010100000000101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110100100111110110111000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111110100000001111010000111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111100000000111101101111101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111110110111110010110001001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111110101101011110111101100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110101011001011111001000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110001001010100001110001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111110010100110000011101001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111101110000010011000011110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111110001110000011110011011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111110101011000110001101101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111101000111100110001111000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111101110110010111100100100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111110110111010000000110010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111111001111010001101000110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111101010101010100110000110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111110110010101101100011110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111110010100110001001111000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel59_Valid_Out)
	);
	Adder_32input add_k59(
		.Data1(Data_Out_Kernel59[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel59[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel59[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel59[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel59[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel59[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel59[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel59[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel59[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel59[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel59[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel59[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel59[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel59[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel59[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel59[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel59[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel59[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel59[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel59[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel59[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel59[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel59[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel59[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel59[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel59[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel59[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel59[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel59[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel59[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel59[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel59[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel59),
		.Data_Out(add_k59_Data_Out),
		.Valid_Out(add_kernel59_Valid_Out)
	);
	Batch_Norm bn_kernel59(
		.Data_A(32'b00111110100011011010111100100100),
		.Data_B(32'b00111110111000100011010001111111),
		.Data_In(add_k59_Data_Out),
		.Valid_In(add_kernel59_Valid_Out),
		.Data_Out(bn59_Data_Out),
		.Valid_Out(bn59_Valid_Out)
	);
	Relu_Core rl_kernel59(
		.Data_In(bn59_Data_Out),
		.Valid_In(bn59_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(rl59_Valid_Out)
	);
//////////KERNEL60//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110100000111011111011000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111110110010001010100010110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110101101101010110000100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111101110000010000000110111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111111010101111100011010110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111111000110111111110001101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111110000100001100111100010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111111000010100111101001010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111101000000100010110110001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111101010010011101010100000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111111011011000011111111011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110101110010111000011001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111110111000000000111010100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111100011101110100011000010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110101001100000010100010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111101111110011011110001100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111110100110001101001010001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110000101110111110010000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111110111010110001110000000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110101111110101010100101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110101101011100100100001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111101110010001011011011010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110011101111010010100100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111110111010000111011010111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111110010110010100111110000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110000001000111111100011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111101100110100011000011001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110000110010010111010101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111110010101011100000111110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110010011010111100101010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111110101101110100101111001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111101010111000001100011100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel60_Valid_Out)
	);
	Adder_32input add_k60(
		.Data1(Data_Out_Kernel60[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel60[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel60[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel60[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel60[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel60[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel60[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel60[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel60[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel60[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel60[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel60[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel60[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel60[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel60[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel60[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel60[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel60[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel60[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel60[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel60[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel60[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel60[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel60[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel60[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel60[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel60[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel60[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel60[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel60[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel60[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel60[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel60),
		.Data_Out(add_k60_Data_Out),
		.Valid_Out(add_kernel60_Valid_Out)
	);
	Batch_Norm bn_kernel60(
		.Data_A(32'b00111110100011110110101111011101),
		.Data_B(32'b00111111000111110000011000110110),
		.Data_In(add_k60_Data_Out),
		.Valid_In(add_kernel60_Valid_Out),
		.Data_Out(bn60_Data_Out),
		.Valid_Out(bn60_Valid_Out)
	);
	Relu_Core rl_kernel60(
		.Data_In(bn60_Data_Out),
		.Valid_In(bn60_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(rl60_Valid_Out)
	);
//////////KERNEL61//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110100111010101110011011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111110100010000110110100010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111011111110000001101010110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111101010110110011000100110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111110011010000010110101101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111111001001110111010011110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111110000010100001001101110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111110100100101000010010001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111110100010001000101010000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110101010000000111001101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111111100010100101001111010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111100101001010000001010111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111111001110000010101000100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111101001111101101001110110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110111111001001010011010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111111000100001111011001100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110010000111010011100100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111110011000001111100010010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111111001001100101100100111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111101101100110111110111101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110100001100010111000010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111110101110110011001100001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110111001001010001110101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111101110000110111101000011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111110110011111100110101100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111111000000110000100010111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111100101110000000100011010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111101111110011110111011101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111101001000110101100111110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110011110101111000111100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111101110101000110111110011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111001110011001101110110010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel61_Valid_Out)
	);
	Adder_32input add_k61(
		.Data1(Data_Out_Kernel61[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel61[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel61[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel61[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel61[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel61[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel61[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel61[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel61[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel61[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel61[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel61[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel61[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel61[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel61[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel61[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel61[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel61[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel61[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel61[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel61[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel61[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel61[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel61[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel61[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel61[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel61[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel61[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel61[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel61[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel61[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel61[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel61),
		.Data_Out(add_k61_Data_Out),
		.Valid_Out(add_kernel61_Valid_Out)
	);
	Batch_Norm bn_kernel61(
		.Data_A(32'b00111110101001110000011100100010),
		.Data_B(32'b10111110100011011010110101011100),
		.Data_In(add_k61_Data_Out),
		.Valid_In(add_kernel61_Valid_Out),
		.Data_Out(bn61_Data_Out),
		.Valid_Out(bn61_Valid_Out)
	);
	Relu_Core rl_kernel61(
		.Data_In(bn61_Data_Out),
		.Valid_In(bn61_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(rl61_Valid_Out)
	);
//////////KERNEL62//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110111010000110011111100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110111000000011001110101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111101111010000001011101011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110100000111001111001000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111101111011101010000110011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110101110001110010001101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111110110100010100000011101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111110111000111110101010011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111110110001101011111001111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110100000000000010001010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110001010101011001000011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111110101111111100001101101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111111001011110100111001101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111110000100000011000011001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110011011101100001111111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111110101000100010101001011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111110000000110011101001100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111110001101101100011010110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111111000010111000010110100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111101100100010110011000001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110100000011010011000000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111110011111011010110011101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111100111101000101111111110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111101101111001110111001100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111111011001111001110110011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111101101001111110111101110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111110101101001000111110011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111110111110010111101010001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111110110111001111111111011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110010000010000001100011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111110111111101110001110110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111101111000101100110001101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel62_Valid_Out)
	);
	Adder_32input add_k62(
		.Data1(Data_Out_Kernel62[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel62[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel62[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel62[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel62[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel62[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel62[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel62[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel62[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel62[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel62[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel62[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel62[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel62[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel62[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel62[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel62[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel62[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel62[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel62[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel62[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel62[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel62[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel62[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel62[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel62[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel62[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel62[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel62[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel62[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel62[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel62[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel62),
		.Data_Out(add_k62_Data_Out),
		.Valid_Out(add_kernel62_Valid_Out)
	);
	Batch_Norm bn_kernel62(
		.Data_A(32'b00111110010001100001000111001111),
		.Data_B(32'b00111110110011110011011111100010),
		.Data_In(add_k62_Data_Out),
		.Valid_In(add_kernel62_Valid_Out),
		.Data_Out(bn62_Data_Out),
		.Valid_Out(bn62_Valid_Out)
	);
	Relu_Core rl_kernel62(
		.Data_In(bn62_Data_Out),
		.Valid_In(bn62_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(rl62_Valid_Out)
	);
//////////KERNEL63//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111110100000011101100100000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111110110111111010100011001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110000111110011000101010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111111000110100110000100111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111111001101111001111010000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110101010000010001111101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111101110100101111011111101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111101100001101001000000111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111110001010100010111001111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111111000001011001111101111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111010110110111010100100001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110010101111100001110011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110101000010111011100000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111110110000001010111000001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110101010111101000001010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111101110000111011011010000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111101010111110011111111100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110100010001000100110100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111101111001101000000111100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111110101011011011101001011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111101110010110010000000101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111110110000011010010110010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110111001100011111011100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111110001001001101100101110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111111001011111000001111011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111101001101100110011001101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110011110100001000111001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111110100010001100110010001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111110011100000101100001001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110110001010111101011100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111110101110010111100010011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111111010101110001100111001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel63_Valid_Out)
	);
	Adder_32input add_k63(
		.Data1(Data_Out_Kernel63[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel63[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel63[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel63[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel63[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel63[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel63[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel63[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel63[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel63[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel63[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel63[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel63[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel63[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel63[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel63[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel63[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel63[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel63[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel63[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel63[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel63[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel63[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel63[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel63[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel63[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel63[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel63[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel63[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel63[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel63[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel63[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel63),
		.Data_Out(add_k63_Data_Out),
		.Valid_Out(add_kernel63_Valid_Out)
	);
	Batch_Norm bn_kernel63(
		.Data_A(32'b00111110101101001100010101000111),
		.Data_B(32'b10111110100000011010000100110000),
		.Data_In(add_k63_Data_Out),
		.Valid_In(add_kernel63_Valid_Out),
		.Data_Out(bn63_Data_Out),
		.Valid_Out(bn63_Valid_Out)
	);
	Relu_Core rl_kernel63(
		.Data_In(bn63_Data_Out),
		.Valid_In(bn63_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(rl63_Valid_Out)
	);
//////////KERNEL64//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110101011010101111110011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111101001100111110110100001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110100101001111000110011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110011011111001100001110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111111000010100101110111011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111110100000101101101101100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111110101101011001011101111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111110011011100001100000000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111010000010100100011011011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110000010001000110011101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111111001010100011010011100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111111001011011110010100000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110111101111100001011001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111110010000010111110100001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110010101001111110111110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111111001000001001001100100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111101000111001110011010111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111010000111000111010011110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111101111001100110111001000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110111010010100111111000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110100011011000000010011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111100010100011110111110000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110101100010001001111001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111110100010111100101010011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111111000100101101100110001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111110100011001001110101001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110000011101110001000000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110001011010001100001101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111111001010000001111111101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111100110110100100100000010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111111000000000010010001000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110100100010010010110011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel64_Valid_Out)
	);
	Adder_32input add_k64(
		.Data1(Data_Out_Kernel64[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel64[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel64[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel64[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel64[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel64[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel64[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel64[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel64[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel64[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel64[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel64[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel64[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel64[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel64[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel64[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel64[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel64[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel64[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel64[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel64[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel64[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel64[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel64[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel64[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel64[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel64[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel64[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel64[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel64[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel64[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel64[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel64),
		.Data_Out(add_k64_Data_Out),
		.Valid_Out(add_kernel64_Valid_Out)
	);
	Batch_Norm bn_kernel64(
		.Data_A(32'b00111110011110010000001100100010),
		.Data_B(32'b10111110000011100000101110111110),
		.Data_In(add_k64_Data_Out),
		.Valid_In(add_kernel64_Valid_Out),
		.Data_Out(bn64_Data_Out),
		.Valid_Out(bn64_Valid_Out)
	);
	Relu_Core rl_kernel64(
		.Data_In(bn64_Data_Out),
		.Valid_In(bn64_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(rl64_Valid_Out)
	);

    
endmodule