module Depthwise_Part1_Separable_8CHANNEL #(
    parameter DATA_WIDHT = 32, 
    parameter IMG_WIDHT = 44,
    parameter IMG_HEIGHT =44
)
(
    input [DATA_WIDHT*16-1:0] Data_In,
    input clk,
    input rst,
    input Valid_In,
    output [DATA_WIDHT*16-1:0] Data_Out,
    output Valid_Out

);
    wire CHANNEL1_Valid_Out, CHANNEL2_Valid_Out, CHANNEL3_Valid_Out, CHANNEL4_Valid_Out, CHANNEL5_Valid_Out, CHANNEL6_Valid_Out, CHANNEL7_Valid_Out, CHANNEL8_Valid_Out, CHANNEL9_Valid_Out, CHANNEL10_Valid_Out, CHANNEL11_Valid_Out, CHANNEL12_Valid_Out, CHANNEL13_Valid_Out, CHANNEL14_Valid_Out, CHANNEL15_Valid_Out, CHANNEL16_Valid_Out;

	assign Valid_Out= CHANNEL1_Valid_Out & CHANNEL2_Valid_Out & CHANNEL3_Valid_Out & CHANNEL4_Valid_Out & CHANNEL5_Valid_Out & CHANNEL6_Valid_Out & CHANNEL7_Valid_Out & CHANNEL8_Valid_Out & CHANNEL9_Valid_Out & CHANNEL10_Valid_Out & CHANNEL11_Valid_Out & CHANNEL12_Valid_Out & CHANNEL13_Valid_Out & CHANNEL14_Valid_Out & CHANNEL15_Valid_Out & CHANNEL16_Valid_Out;


    	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL1 (
			.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
			.Kerne0(32'b10111110001110101011000010100010),
			.Kerne1(32'b10111111011011101110011001110111),
			.Kerne2(32'b10111110110010000000000011011001),
			.Kerne3(32'b00111110101001101110000001111000),
			.Kerne4(32'b10111111000110110100001110011001),
			.Kerne5(32'b00111101001011110111100000111011),
			.Kerne6(32'b10111101100100000100010111111011),
			.Kerne7(32'b00111101110100001100111111000101),
			.Kerne8(32'b00111110011111100110001011010010),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT-1:0]),
			.Valid_Out(CHANNEL1_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL2 (
			.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
			.Kerne0(32'b10111111001000000000111010100111),
			.Kerne1(32'b10111110101011011001101101011110),
			.Kerne2(32'b10111110111100111100001011011010),
			.Kerne3(32'b00111110011110011101100110110001),
			.Kerne4(32'b00111110011110101100010000100010),
			.Kerne5(32'b00111110100110111000101010000011),
			.Kerne6(32'b00111111001110011110110000011110),
			.Kerne7(32'b00111110110011111101100100010110),
			.Kerne8(32'b00111110110010111100001011010001),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*2-1:DATA_WIDHT*1]),
			.Valid_Out(CHANNEL2_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL3 (
			.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
			.Kerne0(32'b10111101111011110010011000110000),
			.Kerne1(32'b10111111010111100101011001000011),
			.Kerne2(32'b00111101001010111100101010100011),
			.Kerne3(32'b10111110110101010110010000101000),
			.Kerne4(32'b00111101101001010111100111010000),
			.Kerne5(32'b10111111000101000101111110011001),
			.Kerne6(32'b00111110101101111001101110010101),
			.Kerne7(32'b00111110100011001011011010001111),
			.Kerne8(32'b10111110100101111011110010011111),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*3-1:DATA_WIDHT*2]),
			.Valid_Out(CHANNEL3_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL4 (
			.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
			.Kerne0(32'b00111110101101101000101111111000),
			.Kerne1(32'b10111111001000010101010001110010),
			.Kerne2(32'b10111110100101111001100001111000),
			.Kerne3(32'b10111110011000101100000001001110),
			.Kerne4(32'b10111110011011100001100001010101),
			.Kerne5(32'b10111110110000110111111110010111),
			.Kerne6(32'b10111110101111001001111001110101),
			.Kerne7(32'b10111100111011010110000011011011),
			.Kerne8(32'b10111110101001111111100101010111),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*4-1:DATA_WIDHT*3]),
			.Valid_Out(CHANNEL4_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL5 (
			.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
			.Kerne0(32'b10111110111111001111110001001110),
			.Kerne1(32'b00111110101010100111010000011101),
			.Kerne2(32'b00111110110010101111000000011011),
			.Kerne3(32'b10111110110011011001110101001001),
			.Kerne4(32'b00111111000110001110001010101011),
			.Kerne5(32'b00111101100100110011110110101000),
			.Kerne6(32'b00111110000011010001100111100110),
			.Kerne7(32'b00111110111100011101100110011100),
			.Kerne8(32'b10111111000001100111010001001000),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*5-1:DATA_WIDHT*4]),
			.Valid_Out(CHANNEL5_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL6 (
			.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
			.Kerne0(32'b10111110100001001000101010001010),
			.Kerne1(32'b00111101101001001010011111100111),
			.Kerne2(32'b00111100001101111010010101110001),
			.Kerne3(32'b10111101110100101100110010100011),
			.Kerne4(32'b10111110100011011000010000011101),
			.Kerne5(32'b00111111000010110110110100100010),
			.Kerne6(32'b00111110001000100111000101001111),
			.Kerne7(32'b00111110101001010110101101100010),
			.Kerne8(32'b00111111010011000010100000111101),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*6-1:DATA_WIDHT*5]),
			.Valid_Out(CHANNEL6_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL7 (
			.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
			.Kerne0(32'b00111101111100011010100001100011),
			.Kerne1(32'b00111110100100101011101011111101),
			.Kerne2(32'b00111110000110101010111001000010),
			.Kerne3(32'b00111101100011111010010101000110),
			.Kerne4(32'b10111101111011010111001011100011),
			.Kerne5(32'b10111110011010110001100110100101),
			.Kerne6(32'b10111110100011101101111011100100),
			.Kerne7(32'b10111111011011010100011110100101),
			.Kerne8(32'b10111110111000011101011001101100),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*7-1:DATA_WIDHT*6]),
			.Valid_Out(CHANNEL7_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL8 (
			.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
			.Kerne0(32'b10111100000111011110110010101001),
			.Kerne1(32'b00111110111010011101111001100100),
			.Kerne2(32'b10111101100100010100010100110101),
			.Kerne3(32'b00111111000110010101001010001011),
			.Kerne4(32'b10111011010000101001110001011001),
			.Kerne5(32'b00111011001110001110110001110001),
			.Kerne6(32'b00111111000011110100111100111100),
			.Kerne7(32'b10111111000000101101100000111110),
			.Kerne8(32'b10111110110101000001001011111100),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*8-1:DATA_WIDHT*7]),
			.Valid_Out(CHANNEL8_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL9 (
			.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
			.Kerne0(32'b10111101001110011010111100100011),
			.Kerne1(32'b00111110101011100000101011000111),
			.Kerne2(32'b10111101110101100101001010000010),
			.Kerne3(32'b00111110111111100000000101110100),
			.Kerne4(32'b10111101101110100101000000111100),
			.Kerne5(32'b00111111000000101010000001111001),
			.Kerne6(32'b00111110000100100101101101110110),
			.Kerne7(32'b10111111000010110101010101001111),
			.Kerne8(32'b10111111001111101110111010001101),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*9-1:DATA_WIDHT*8]),
			.Valid_Out(CHANNEL9_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL10 (
			.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
			.Kerne0(32'b00111110111001010000111110000010),
			.Kerne1(32'b00111110100010110000001110000101),
			.Kerne2(32'b00111110001011100100111011110001),
			.Kerne3(32'b00111111000001111111101111010001),
			.Kerne4(32'b00111110111011000011010010000001),
			.Kerne5(32'b00111110100110111110110110000101),
			.Kerne6(32'b00111110101010110101000101110100),
			.Kerne7(32'b10111110011100000100000100011100),
			.Kerne8(32'b00111110111000000101000110101011),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*10-1:DATA_WIDHT*9]),
			.Valid_Out(CHANNEL10_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL11 (
			.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
			.Kerne0(32'b10111110110100111001111001111111),
			.Kerne1(32'b00111110100100011111101100010110),
			.Kerne2(32'b00111110000011100100010101001010),
			.Kerne3(32'b10111111010000100011110010100010),
			.Kerne4(32'b10111110011011001001000010000101),
			.Kerne5(32'b00111110101010101000101111110001),
			.Kerne6(32'b10111110110010011010111001011111),
			.Kerne7(32'b00111101011100001111100010111011),
			.Kerne8(32'b00111111000101111000110000000010),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*11-1:DATA_WIDHT*10]),
			.Valid_Out(CHANNEL11_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL12 (
			.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
			.Kerne0(32'b00111110000101011100101000111110),
			.Kerne1(32'b00111111001111010100010101101110),
			.Kerne2(32'b10111101001000110011101001101101),
			.Kerne3(32'b00111111000001000100111011010001),
			.Kerne4(32'b00111111001100001110000001010100),
			.Kerne5(32'b10111110101010100001100000011010),
			.Kerne6(32'b10111101010010100110110001010001),
			.Kerne7(32'b00111101000110011001001001100011),
			.Kerne8(32'b10111010100001011100101100110010),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*12-1:DATA_WIDHT*11]),
			.Valid_Out(CHANNEL12_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL13 (
			.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
			.Kerne0(32'b10111110110110000100001010010010),
			.Kerne1(32'b00111110000010011010111110101100),
			.Kerne2(32'b10111111010011100010110000010001),
			.Kerne3(32'b00111101101011111001111000011100),
			.Kerne4(32'b10111101011101111011111110000000),
			.Kerne5(32'b00111110111001111000100101010010),
			.Kerne6(32'b00111110100111001001010111010001),
			.Kerne7(32'b10111110101100110010110101001111),
			.Kerne8(32'b00111110110100110001010011011100),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*13-1:DATA_WIDHT*12]),
			.Valid_Out(CHANNEL13_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL14 (
			.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
			.Kerne0(32'b00111101100010011111010111101011),
			.Kerne1(32'b00111111011011100101000010110010),
			.Kerne2(32'b00111110001111000110111111011100),
			.Kerne3(32'b10111110000000010111000101000101),
			.Kerne4(32'b00111110101110011000101100100100),
			.Kerne5(32'b00111111000110010101011001111111),
			.Kerne6(32'b00111110011001101110101110110011),
			.Kerne7(32'b00111101001010110000011010110100),
			.Kerne8(32'b00111110101000110011110000000000),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*14-1:DATA_WIDHT*13]),
			.Valid_Out(CHANNEL14_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL15 (
			.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
			.Kerne0(32'b10111101110010011011101100011101),
			.Kerne1(32'b00111111011100001001011100001000),
			.Kerne2(32'b10111110000011000010010001111011),
			.Kerne3(32'b00111100001000100010111010100000),
			.Kerne4(32'b00111110011110101101001001111111),
			.Kerne5(32'b10111110100101111001010010110100),
			.Kerne6(32'b10111110101010011110010111101011),
			.Kerne7(32'b10111110011111011010001111000100),
			.Kerne8(32'b10111110101111110101100110111000),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*15-1:DATA_WIDHT*14]),
			.Valid_Out(CHANNEL15_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL16 (
			.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
			.Kerne0(32'b00111110011011111110111110000001),
			.Kerne1(32'b00111110011101000001010001010010),
			.Kerne2(32'b00111110110000000101100011110011),
			.Kerne3(32'b00111110101100101110111011001111),
			.Kerne4(32'b10111101000101111111000101010100),
			.Kerne5(32'b00111110101010110110011100001001),
			.Kerne6(32'b00111110110011110111011101101000),
			.Kerne7(32'b10111101001111100111011000010010),
			.Kerne8(32'b00111111010000101101011111110100),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*16-1:DATA_WIDHT*15]),
			.Valid_Out(CHANNEL16_Valid_Out)
		);

endmodule