// module Adder_GAVG #(
//     parameter DATA_WIDHT = 32,
//     parameter SUM = 20;
// ) (
//     input [31:0] Data_In,
//     input Valid_In,
//     output [31:0] Data_Out,
//     output Valid_Out
// );
//     reg[31:0] Counter = 0;
//     always @() begin
        
//     end
//     always @(Valid_In or Data_In) begin
    
//     end
    
// endmodule