module Depthwise_Part3_Separable_64CHANNEL_Layer5 #(
    parameter DATA_WIDHT = 32, 
    parameter IMG_WIDHT = 44,
    parameter IMG_HEIGHT =44
)
(
    input [DATA_WIDHT*64-1:0] Data_In,
    input clk,
    input rst,
    input Valid_In,
    output [DATA_WIDHT*64-1:0] Data_Out,
    output Valid_Out

);
	wire[DATA_WIDHT*64-1:0] Data_Out_Kernel1, Data_Out_Kernel2, Data_Out_Kernel3, Data_Out_Kernel4, Data_Out_Kernel5, Data_Out_Kernel6, Data_Out_Kernel7, Data_Out_Kernel8, Data_Out_Kernel9, Data_Out_Kernel10, Data_Out_Kernel11, Data_Out_Kernel12, Data_Out_Kernel13, Data_Out_Kernel14, Data_Out_Kernel15, Data_Out_Kernel16, Data_Out_Kernel17, Data_Out_Kernel18, Data_Out_Kernel19, Data_Out_Kernel20, Data_Out_Kernel21, Data_Out_Kernel22, Data_Out_Kernel23, Data_Out_Kernel24, Data_Out_Kernel25, Data_Out_Kernel26, Data_Out_Kernel27, Data_Out_Kernel28, Data_Out_Kernel29, Data_Out_Kernel30, Data_Out_Kernel31, Data_Out_Kernel32, Data_Out_Kernel33, Data_Out_Kernel34, Data_Out_Kernel35, Data_Out_Kernel36, Data_Out_Kernel37, Data_Out_Kernel38, Data_Out_Kernel39, Data_Out_Kernel40, Data_Out_Kernel41, Data_Out_Kernel42, Data_Out_Kernel43, Data_Out_Kernel44, Data_Out_Kernel45, Data_Out_Kernel46, Data_Out_Kernel47, Data_Out_Kernel48, Data_Out_Kernel49, Data_Out_Kernel50, Data_Out_Kernel51, Data_Out_Kernel52, Data_Out_Kernel53, Data_Out_Kernel54, Data_Out_Kernel55, Data_Out_Kernel56, Data_Out_Kernel57, Data_Out_Kernel58, Data_Out_Kernel59, Data_Out_Kernel60, Data_Out_Kernel61, Data_Out_Kernel62, Data_Out_Kernel63, Data_Out_Kernel64;
	
	wire[31:0] add_k1_Data_Out, add_k2_Data_Out, add_k3_Data_Out, add_k4_Data_Out, add_k5_Data_Out, add_k6_Data_Out, add_k7_Data_Out, add_k8_Data_Out, add_k9_Data_Out, add_k10_Data_Out, add_k11_Data_Out, add_k12_Data_Out, add_k13_Data_Out, add_k14_Data_Out, add_k15_Data_Out, add_k16_Data_Out, add_k17_Data_Out, add_k18_Data_Out, add_k19_Data_Out, add_k20_Data_Out, add_k21_Data_Out, add_k22_Data_Out, add_k23_Data_Out, add_k24_Data_Out, add_k25_Data_Out, add_k26_Data_Out, add_k27_Data_Out, add_k28_Data_Out, add_k29_Data_Out, add_k30_Data_Out, add_k31_Data_Out, add_k32_Data_Out, add_k33_Data_Out, add_k34_Data_Out, add_k35_Data_Out, add_k36_Data_Out, add_k37_Data_Out, add_k38_Data_Out, add_k39_Data_Out, add_k40_Data_Out, add_k41_Data_Out, add_k42_Data_Out, add_k43_Data_Out, add_k44_Data_Out, add_k45_Data_Out, add_k46_Data_Out, add_k47_Data_Out, add_k48_Data_Out, add_k49_Data_Out, add_k50_Data_Out, add_k51_Data_Out, add_k52_Data_Out, add_k53_Data_Out, add_k54_Data_Out, add_k55_Data_Out, add_k56_Data_Out, add_k57_Data_Out, add_k58_Data_Out, add_k59_Data_Out, add_k60_Data_Out, add_k61_Data_Out, add_k62_Data_Out, add_k63_Data_Out, add_k64_Data_Out;

	wire add_kernel1_Valid_Out, add_kernel2_Valid_Out, add_kernel3_Valid_Out, add_kernel4_Valid_Out, add_kernel5_Valid_Out, add_kernel6_Valid_Out, add_kernel7_Valid_Out, add_kernel8_Valid_Out, add_kernel9_Valid_Out, add_kernel10_Valid_Out, add_kernel11_Valid_Out, add_kernel12_Valid_Out, add_kernel13_Valid_Out, add_kernel14_Valid_Out, add_kernel15_Valid_Out, add_kernel16_Valid_Out, add_kernel17_Valid_Out, add_kernel18_Valid_Out, add_kernel19_Valid_Out, add_kernel20_Valid_Out, add_kernel21_Valid_Out, add_kernel22_Valid_Out, add_kernel23_Valid_Out, add_kernel24_Valid_Out, add_kernel25_Valid_Out, add_kernel26_Valid_Out, add_kernel27_Valid_Out, add_kernel28_Valid_Out, add_kernel29_Valid_Out, add_kernel30_Valid_Out, add_kernel31_Valid_Out, add_kernel32_Valid_Out, add_kernel33_Valid_Out, add_kernel34_Valid_Out, add_kernel35_Valid_Out, add_kernel36_Valid_Out, add_kernel37_Valid_Out, add_kernel38_Valid_Out, add_kernel39_Valid_Out, add_kernel40_Valid_Out, add_kernel41_Valid_Out, add_kernel42_Valid_Out, add_kernel43_Valid_Out, add_kernel44_Valid_Out, add_kernel45_Valid_Out, add_kernel46_Valid_Out, add_kernel47_Valid_Out, add_kernel48_Valid_Out, add_kernel49_Valid_Out, add_kernel50_Valid_Out, add_kernel51_Valid_Out, add_kernel52_Valid_Out, add_kernel53_Valid_Out, add_kernel54_Valid_Out, add_kernel55_Valid_Out, add_kernel56_Valid_Out, add_kernel57_Valid_Out, add_kernel58_Valid_Out, add_kernel59_Valid_Out, add_kernel60_Valid_Out, add_kernel61_Valid_Out, add_kernel62_Valid_Out, add_kernel63_Valid_Out, add_kernel64_Valid_Out;

	wire channel1_Kernel1_Valid_Out, channel2_Kernel1_Valid_Out, channel3_Kernel1_Valid_Out, channel4_Kernel1_Valid_Out, channel5_Kernel1_Valid_Out, channel6_Kernel1_Valid_Out, channel7_Kernel1_Valid_Out, channel8_Kernel1_Valid_Out, channel9_Kernel1_Valid_Out, channel10_Kernel1_Valid_Out, channel11_Kernel1_Valid_Out, channel12_Kernel1_Valid_Out, channel13_Kernel1_Valid_Out, channel14_Kernel1_Valid_Out, channel15_Kernel1_Valid_Out, channel16_Kernel1_Valid_Out, channel17_Kernel1_Valid_Out, channel18_Kernel1_Valid_Out, channel19_Kernel1_Valid_Out, channel20_Kernel1_Valid_Out, channel21_Kernel1_Valid_Out, channel22_Kernel1_Valid_Out, channel23_Kernel1_Valid_Out, channel24_Kernel1_Valid_Out, channel25_Kernel1_Valid_Out, channel26_Kernel1_Valid_Out, channel27_Kernel1_Valid_Out, channel28_Kernel1_Valid_Out, channel29_Kernel1_Valid_Out, channel30_Kernel1_Valid_Out, channel31_Kernel1_Valid_Out, channel32_Kernel1_Valid_Out, channel33_Kernel1_Valid_Out, channel34_Kernel1_Valid_Out, channel35_Kernel1_Valid_Out, channel36_Kernel1_Valid_Out, channel37_Kernel1_Valid_Out, channel38_Kernel1_Valid_Out, channel39_Kernel1_Valid_Out, channel40_Kernel1_Valid_Out, channel41_Kernel1_Valid_Out, channel42_Kernel1_Valid_Out, channel43_Kernel1_Valid_Out, channel44_Kernel1_Valid_Out, channel45_Kernel1_Valid_Out, channel46_Kernel1_Valid_Out, channel47_Kernel1_Valid_Out, channel48_Kernel1_Valid_Out, channel49_Kernel1_Valid_Out, channel50_Kernel1_Valid_Out, channel51_Kernel1_Valid_Out, channel52_Kernel1_Valid_Out, channel53_Kernel1_Valid_Out, channel54_Kernel1_Valid_Out, channel55_Kernel1_Valid_Out, channel56_Kernel1_Valid_Out, channel57_Kernel1_Valid_Out, channel58_Kernel1_Valid_Out, channel59_Kernel1_Valid_Out, channel60_Kernel1_Valid_Out, channel61_Kernel1_Valid_Out, channel62_Kernel1_Valid_Out, channel63_Kernel1_Valid_Out, channel64_Kernel1_Valid_Out;

	assign add_kernel1=channel1_Kernel1_Valid_Out & channel2_Kernel1_Valid_Out & channel3_Kernel1_Valid_Out & channel4_Kernel1_Valid_Out & channel5_Kernel1_Valid_Out & channel6_Kernel1_Valid_Out & channel7_Kernel1_Valid_Out & channel8_Kernel1_Valid_Out & channel9_Kernel1_Valid_Out & channel10_Kernel1_Valid_Out & channel11_Kernel1_Valid_Out & channel12_Kernel1_Valid_Out & channel13_Kernel1_Valid_Out & channel14_Kernel1_Valid_Out & channel15_Kernel1_Valid_Out & channel16_Kernel1_Valid_Out & channel17_Kernel1_Valid_Out & channel18_Kernel1_Valid_Out & channel19_Kernel1_Valid_Out & channel20_Kernel1_Valid_Out & channel21_Kernel1_Valid_Out & channel22_Kernel1_Valid_Out & channel23_Kernel1_Valid_Out & channel24_Kernel1_Valid_Out & channel25_Kernel1_Valid_Out & channel26_Kernel1_Valid_Out & channel27_Kernel1_Valid_Out & channel28_Kernel1_Valid_Out & channel29_Kernel1_Valid_Out & channel30_Kernel1_Valid_Out & channel31_Kernel1_Valid_Out & channel32_Kernel1_Valid_Out & channel33_Kernel1_Valid_Out & channel34_Kernel1_Valid_Out & channel35_Kernel1_Valid_Out & channel36_Kernel1_Valid_Out & channel37_Kernel1_Valid_Out & channel38_Kernel1_Valid_Out & channel39_Kernel1_Valid_Out & channel40_Kernel1_Valid_Out & channel41_Kernel1_Valid_Out & channel42_Kernel1_Valid_Out & channel43_Kernel1_Valid_Out & channel44_Kernel1_Valid_Out & channel45_Kernel1_Valid_Out & channel46_Kernel1_Valid_Out & channel47_Kernel1_Valid_Out & channel48_Kernel1_Valid_Out & channel49_Kernel1_Valid_Out & channel50_Kernel1_Valid_Out & channel51_Kernel1_Valid_Out & channel52_Kernel1_Valid_Out & channel53_Kernel1_Valid_Out & channel54_Kernel1_Valid_Out & channel55_Kernel1_Valid_Out & channel56_Kernel1_Valid_Out & channel57_Kernel1_Valid_Out & channel58_Kernel1_Valid_Out & channel59_Kernel1_Valid_Out & channel60_Kernel1_Valid_Out & channel61_Kernel1_Valid_Out & channel62_Kernel1_Valid_Out & channel63_Kernel1_Valid_Out & channel64_Kernel1_Valid_Out;

	wire channel1_Kernel2_Valid_Out, channel2_Kernel2_Valid_Out, channel3_Kernel2_Valid_Out, channel4_Kernel2_Valid_Out, channel5_Kernel2_Valid_Out, channel6_Kernel2_Valid_Out, channel7_Kernel2_Valid_Out, channel8_Kernel2_Valid_Out, channel9_Kernel2_Valid_Out, channel10_Kernel2_Valid_Out, channel11_Kernel2_Valid_Out, channel12_Kernel2_Valid_Out, channel13_Kernel2_Valid_Out, channel14_Kernel2_Valid_Out, channel15_Kernel2_Valid_Out, channel16_Kernel2_Valid_Out, channel17_Kernel2_Valid_Out, channel18_Kernel2_Valid_Out, channel19_Kernel2_Valid_Out, channel20_Kernel2_Valid_Out, channel21_Kernel2_Valid_Out, channel22_Kernel2_Valid_Out, channel23_Kernel2_Valid_Out, channel24_Kernel2_Valid_Out, channel25_Kernel2_Valid_Out, channel26_Kernel2_Valid_Out, channel27_Kernel2_Valid_Out, channel28_Kernel2_Valid_Out, channel29_Kernel2_Valid_Out, channel30_Kernel2_Valid_Out, channel31_Kernel2_Valid_Out, channel32_Kernel2_Valid_Out, channel33_Kernel2_Valid_Out, channel34_Kernel2_Valid_Out, channel35_Kernel2_Valid_Out, channel36_Kernel2_Valid_Out, channel37_Kernel2_Valid_Out, channel38_Kernel2_Valid_Out, channel39_Kernel2_Valid_Out, channel40_Kernel2_Valid_Out, channel41_Kernel2_Valid_Out, channel42_Kernel2_Valid_Out, channel43_Kernel2_Valid_Out, channel44_Kernel2_Valid_Out, channel45_Kernel2_Valid_Out, channel46_Kernel2_Valid_Out, channel47_Kernel2_Valid_Out, channel48_Kernel2_Valid_Out, channel49_Kernel2_Valid_Out, channel50_Kernel2_Valid_Out, channel51_Kernel2_Valid_Out, channel52_Kernel2_Valid_Out, channel53_Kernel2_Valid_Out, channel54_Kernel2_Valid_Out, channel55_Kernel2_Valid_Out, channel56_Kernel2_Valid_Out, channel57_Kernel2_Valid_Out, channel58_Kernel2_Valid_Out, channel59_Kernel2_Valid_Out, channel60_Kernel2_Valid_Out, channel61_Kernel2_Valid_Out, channel62_Kernel2_Valid_Out, channel63_Kernel2_Valid_Out, channel64_Kernel2_Valid_Out;

	assign add_kernel2=channel1_Kernel2_Valid_Out & channel2_Kernel2_Valid_Out & channel3_Kernel2_Valid_Out & channel4_Kernel2_Valid_Out & channel5_Kernel2_Valid_Out & channel6_Kernel2_Valid_Out & channel7_Kernel2_Valid_Out & channel8_Kernel2_Valid_Out & channel9_Kernel2_Valid_Out & channel10_Kernel2_Valid_Out & channel11_Kernel2_Valid_Out & channel12_Kernel2_Valid_Out & channel13_Kernel2_Valid_Out & channel14_Kernel2_Valid_Out & channel15_Kernel2_Valid_Out & channel16_Kernel2_Valid_Out & channel17_Kernel2_Valid_Out & channel18_Kernel2_Valid_Out & channel19_Kernel2_Valid_Out & channel20_Kernel2_Valid_Out & channel21_Kernel2_Valid_Out & channel22_Kernel2_Valid_Out & channel23_Kernel2_Valid_Out & channel24_Kernel2_Valid_Out & channel25_Kernel2_Valid_Out & channel26_Kernel2_Valid_Out & channel27_Kernel2_Valid_Out & channel28_Kernel2_Valid_Out & channel29_Kernel2_Valid_Out & channel30_Kernel2_Valid_Out & channel31_Kernel2_Valid_Out & channel32_Kernel2_Valid_Out & channel33_Kernel2_Valid_Out & channel34_Kernel2_Valid_Out & channel35_Kernel2_Valid_Out & channel36_Kernel2_Valid_Out & channel37_Kernel2_Valid_Out & channel38_Kernel2_Valid_Out & channel39_Kernel2_Valid_Out & channel40_Kernel2_Valid_Out & channel41_Kernel2_Valid_Out & channel42_Kernel2_Valid_Out & channel43_Kernel2_Valid_Out & channel44_Kernel2_Valid_Out & channel45_Kernel2_Valid_Out & channel46_Kernel2_Valid_Out & channel47_Kernel2_Valid_Out & channel48_Kernel2_Valid_Out & channel49_Kernel2_Valid_Out & channel50_Kernel2_Valid_Out & channel51_Kernel2_Valid_Out & channel52_Kernel2_Valid_Out & channel53_Kernel2_Valid_Out & channel54_Kernel2_Valid_Out & channel55_Kernel2_Valid_Out & channel56_Kernel2_Valid_Out & channel57_Kernel2_Valid_Out & channel58_Kernel2_Valid_Out & channel59_Kernel2_Valid_Out & channel60_Kernel2_Valid_Out & channel61_Kernel2_Valid_Out & channel62_Kernel2_Valid_Out & channel63_Kernel2_Valid_Out & channel64_Kernel2_Valid_Out;

	wire channel1_Kernel3_Valid_Out, channel2_Kernel3_Valid_Out, channel3_Kernel3_Valid_Out, channel4_Kernel3_Valid_Out, channel5_Kernel3_Valid_Out, channel6_Kernel3_Valid_Out, channel7_Kernel3_Valid_Out, channel8_Kernel3_Valid_Out, channel9_Kernel3_Valid_Out, channel10_Kernel3_Valid_Out, channel11_Kernel3_Valid_Out, channel12_Kernel3_Valid_Out, channel13_Kernel3_Valid_Out, channel14_Kernel3_Valid_Out, channel15_Kernel3_Valid_Out, channel16_Kernel3_Valid_Out, channel17_Kernel3_Valid_Out, channel18_Kernel3_Valid_Out, channel19_Kernel3_Valid_Out, channel20_Kernel3_Valid_Out, channel21_Kernel3_Valid_Out, channel22_Kernel3_Valid_Out, channel23_Kernel3_Valid_Out, channel24_Kernel3_Valid_Out, channel25_Kernel3_Valid_Out, channel26_Kernel3_Valid_Out, channel27_Kernel3_Valid_Out, channel28_Kernel3_Valid_Out, channel29_Kernel3_Valid_Out, channel30_Kernel3_Valid_Out, channel31_Kernel3_Valid_Out, channel32_Kernel3_Valid_Out, channel33_Kernel3_Valid_Out, channel34_Kernel3_Valid_Out, channel35_Kernel3_Valid_Out, channel36_Kernel3_Valid_Out, channel37_Kernel3_Valid_Out, channel38_Kernel3_Valid_Out, channel39_Kernel3_Valid_Out, channel40_Kernel3_Valid_Out, channel41_Kernel3_Valid_Out, channel42_Kernel3_Valid_Out, channel43_Kernel3_Valid_Out, channel44_Kernel3_Valid_Out, channel45_Kernel3_Valid_Out, channel46_Kernel3_Valid_Out, channel47_Kernel3_Valid_Out, channel48_Kernel3_Valid_Out, channel49_Kernel3_Valid_Out, channel50_Kernel3_Valid_Out, channel51_Kernel3_Valid_Out, channel52_Kernel3_Valid_Out, channel53_Kernel3_Valid_Out, channel54_Kernel3_Valid_Out, channel55_Kernel3_Valid_Out, channel56_Kernel3_Valid_Out, channel57_Kernel3_Valid_Out, channel58_Kernel3_Valid_Out, channel59_Kernel3_Valid_Out, channel60_Kernel3_Valid_Out, channel61_Kernel3_Valid_Out, channel62_Kernel3_Valid_Out, channel63_Kernel3_Valid_Out, channel64_Kernel3_Valid_Out;

	assign add_kernel3=channel1_Kernel3_Valid_Out & channel2_Kernel3_Valid_Out & channel3_Kernel3_Valid_Out & channel4_Kernel3_Valid_Out & channel5_Kernel3_Valid_Out & channel6_Kernel3_Valid_Out & channel7_Kernel3_Valid_Out & channel8_Kernel3_Valid_Out & channel9_Kernel3_Valid_Out & channel10_Kernel3_Valid_Out & channel11_Kernel3_Valid_Out & channel12_Kernel3_Valid_Out & channel13_Kernel3_Valid_Out & channel14_Kernel3_Valid_Out & channel15_Kernel3_Valid_Out & channel16_Kernel3_Valid_Out & channel17_Kernel3_Valid_Out & channel18_Kernel3_Valid_Out & channel19_Kernel3_Valid_Out & channel20_Kernel3_Valid_Out & channel21_Kernel3_Valid_Out & channel22_Kernel3_Valid_Out & channel23_Kernel3_Valid_Out & channel24_Kernel3_Valid_Out & channel25_Kernel3_Valid_Out & channel26_Kernel3_Valid_Out & channel27_Kernel3_Valid_Out & channel28_Kernel3_Valid_Out & channel29_Kernel3_Valid_Out & channel30_Kernel3_Valid_Out & channel31_Kernel3_Valid_Out & channel32_Kernel3_Valid_Out & channel33_Kernel3_Valid_Out & channel34_Kernel3_Valid_Out & channel35_Kernel3_Valid_Out & channel36_Kernel3_Valid_Out & channel37_Kernel3_Valid_Out & channel38_Kernel3_Valid_Out & channel39_Kernel3_Valid_Out & channel40_Kernel3_Valid_Out & channel41_Kernel3_Valid_Out & channel42_Kernel3_Valid_Out & channel43_Kernel3_Valid_Out & channel44_Kernel3_Valid_Out & channel45_Kernel3_Valid_Out & channel46_Kernel3_Valid_Out & channel47_Kernel3_Valid_Out & channel48_Kernel3_Valid_Out & channel49_Kernel3_Valid_Out & channel50_Kernel3_Valid_Out & channel51_Kernel3_Valid_Out & channel52_Kernel3_Valid_Out & channel53_Kernel3_Valid_Out & channel54_Kernel3_Valid_Out & channel55_Kernel3_Valid_Out & channel56_Kernel3_Valid_Out & channel57_Kernel3_Valid_Out & channel58_Kernel3_Valid_Out & channel59_Kernel3_Valid_Out & channel60_Kernel3_Valid_Out & channel61_Kernel3_Valid_Out & channel62_Kernel3_Valid_Out & channel63_Kernel3_Valid_Out & channel64_Kernel3_Valid_Out;

	wire channel1_Kernel4_Valid_Out, channel2_Kernel4_Valid_Out, channel3_Kernel4_Valid_Out, channel4_Kernel4_Valid_Out, channel5_Kernel4_Valid_Out, channel6_Kernel4_Valid_Out, channel7_Kernel4_Valid_Out, channel8_Kernel4_Valid_Out, channel9_Kernel4_Valid_Out, channel10_Kernel4_Valid_Out, channel11_Kernel4_Valid_Out, channel12_Kernel4_Valid_Out, channel13_Kernel4_Valid_Out, channel14_Kernel4_Valid_Out, channel15_Kernel4_Valid_Out, channel16_Kernel4_Valid_Out, channel17_Kernel4_Valid_Out, channel18_Kernel4_Valid_Out, channel19_Kernel4_Valid_Out, channel20_Kernel4_Valid_Out, channel21_Kernel4_Valid_Out, channel22_Kernel4_Valid_Out, channel23_Kernel4_Valid_Out, channel24_Kernel4_Valid_Out, channel25_Kernel4_Valid_Out, channel26_Kernel4_Valid_Out, channel27_Kernel4_Valid_Out, channel28_Kernel4_Valid_Out, channel29_Kernel4_Valid_Out, channel30_Kernel4_Valid_Out, channel31_Kernel4_Valid_Out, channel32_Kernel4_Valid_Out, channel33_Kernel4_Valid_Out, channel34_Kernel4_Valid_Out, channel35_Kernel4_Valid_Out, channel36_Kernel4_Valid_Out, channel37_Kernel4_Valid_Out, channel38_Kernel4_Valid_Out, channel39_Kernel4_Valid_Out, channel40_Kernel4_Valid_Out, channel41_Kernel4_Valid_Out, channel42_Kernel4_Valid_Out, channel43_Kernel4_Valid_Out, channel44_Kernel4_Valid_Out, channel45_Kernel4_Valid_Out, channel46_Kernel4_Valid_Out, channel47_Kernel4_Valid_Out, channel48_Kernel4_Valid_Out, channel49_Kernel4_Valid_Out, channel50_Kernel4_Valid_Out, channel51_Kernel4_Valid_Out, channel52_Kernel4_Valid_Out, channel53_Kernel4_Valid_Out, channel54_Kernel4_Valid_Out, channel55_Kernel4_Valid_Out, channel56_Kernel4_Valid_Out, channel57_Kernel4_Valid_Out, channel58_Kernel4_Valid_Out, channel59_Kernel4_Valid_Out, channel60_Kernel4_Valid_Out, channel61_Kernel4_Valid_Out, channel62_Kernel4_Valid_Out, channel63_Kernel4_Valid_Out, channel64_Kernel4_Valid_Out;

	assign add_kernel4=channel1_Kernel4_Valid_Out & channel2_Kernel4_Valid_Out & channel3_Kernel4_Valid_Out & channel4_Kernel4_Valid_Out & channel5_Kernel4_Valid_Out & channel6_Kernel4_Valid_Out & channel7_Kernel4_Valid_Out & channel8_Kernel4_Valid_Out & channel9_Kernel4_Valid_Out & channel10_Kernel4_Valid_Out & channel11_Kernel4_Valid_Out & channel12_Kernel4_Valid_Out & channel13_Kernel4_Valid_Out & channel14_Kernel4_Valid_Out & channel15_Kernel4_Valid_Out & channel16_Kernel4_Valid_Out & channel17_Kernel4_Valid_Out & channel18_Kernel4_Valid_Out & channel19_Kernel4_Valid_Out & channel20_Kernel4_Valid_Out & channel21_Kernel4_Valid_Out & channel22_Kernel4_Valid_Out & channel23_Kernel4_Valid_Out & channel24_Kernel4_Valid_Out & channel25_Kernel4_Valid_Out & channel26_Kernel4_Valid_Out & channel27_Kernel4_Valid_Out & channel28_Kernel4_Valid_Out & channel29_Kernel4_Valid_Out & channel30_Kernel4_Valid_Out & channel31_Kernel4_Valid_Out & channel32_Kernel4_Valid_Out & channel33_Kernel4_Valid_Out & channel34_Kernel4_Valid_Out & channel35_Kernel4_Valid_Out & channel36_Kernel4_Valid_Out & channel37_Kernel4_Valid_Out & channel38_Kernel4_Valid_Out & channel39_Kernel4_Valid_Out & channel40_Kernel4_Valid_Out & channel41_Kernel4_Valid_Out & channel42_Kernel4_Valid_Out & channel43_Kernel4_Valid_Out & channel44_Kernel4_Valid_Out & channel45_Kernel4_Valid_Out & channel46_Kernel4_Valid_Out & channel47_Kernel4_Valid_Out & channel48_Kernel4_Valid_Out & channel49_Kernel4_Valid_Out & channel50_Kernel4_Valid_Out & channel51_Kernel4_Valid_Out & channel52_Kernel4_Valid_Out & channel53_Kernel4_Valid_Out & channel54_Kernel4_Valid_Out & channel55_Kernel4_Valid_Out & channel56_Kernel4_Valid_Out & channel57_Kernel4_Valid_Out & channel58_Kernel4_Valid_Out & channel59_Kernel4_Valid_Out & channel60_Kernel4_Valid_Out & channel61_Kernel4_Valid_Out & channel62_Kernel4_Valid_Out & channel63_Kernel4_Valid_Out & channel64_Kernel4_Valid_Out;

	wire channel1_Kernel5_Valid_Out, channel2_Kernel5_Valid_Out, channel3_Kernel5_Valid_Out, channel4_Kernel5_Valid_Out, channel5_Kernel5_Valid_Out, channel6_Kernel5_Valid_Out, channel7_Kernel5_Valid_Out, channel8_Kernel5_Valid_Out, channel9_Kernel5_Valid_Out, channel10_Kernel5_Valid_Out, channel11_Kernel5_Valid_Out, channel12_Kernel5_Valid_Out, channel13_Kernel5_Valid_Out, channel14_Kernel5_Valid_Out, channel15_Kernel5_Valid_Out, channel16_Kernel5_Valid_Out, channel17_Kernel5_Valid_Out, channel18_Kernel5_Valid_Out, channel19_Kernel5_Valid_Out, channel20_Kernel5_Valid_Out, channel21_Kernel5_Valid_Out, channel22_Kernel5_Valid_Out, channel23_Kernel5_Valid_Out, channel24_Kernel5_Valid_Out, channel25_Kernel5_Valid_Out, channel26_Kernel5_Valid_Out, channel27_Kernel5_Valid_Out, channel28_Kernel5_Valid_Out, channel29_Kernel5_Valid_Out, channel30_Kernel5_Valid_Out, channel31_Kernel5_Valid_Out, channel32_Kernel5_Valid_Out, channel33_Kernel5_Valid_Out, channel34_Kernel5_Valid_Out, channel35_Kernel5_Valid_Out, channel36_Kernel5_Valid_Out, channel37_Kernel5_Valid_Out, channel38_Kernel5_Valid_Out, channel39_Kernel5_Valid_Out, channel40_Kernel5_Valid_Out, channel41_Kernel5_Valid_Out, channel42_Kernel5_Valid_Out, channel43_Kernel5_Valid_Out, channel44_Kernel5_Valid_Out, channel45_Kernel5_Valid_Out, channel46_Kernel5_Valid_Out, channel47_Kernel5_Valid_Out, channel48_Kernel5_Valid_Out, channel49_Kernel5_Valid_Out, channel50_Kernel5_Valid_Out, channel51_Kernel5_Valid_Out, channel52_Kernel5_Valid_Out, channel53_Kernel5_Valid_Out, channel54_Kernel5_Valid_Out, channel55_Kernel5_Valid_Out, channel56_Kernel5_Valid_Out, channel57_Kernel5_Valid_Out, channel58_Kernel5_Valid_Out, channel59_Kernel5_Valid_Out, channel60_Kernel5_Valid_Out, channel61_Kernel5_Valid_Out, channel62_Kernel5_Valid_Out, channel63_Kernel5_Valid_Out, channel64_Kernel5_Valid_Out;

	assign add_kernel5=channel1_Kernel5_Valid_Out & channel2_Kernel5_Valid_Out & channel3_Kernel5_Valid_Out & channel4_Kernel5_Valid_Out & channel5_Kernel5_Valid_Out & channel6_Kernel5_Valid_Out & channel7_Kernel5_Valid_Out & channel8_Kernel5_Valid_Out & channel9_Kernel5_Valid_Out & channel10_Kernel5_Valid_Out & channel11_Kernel5_Valid_Out & channel12_Kernel5_Valid_Out & channel13_Kernel5_Valid_Out & channel14_Kernel5_Valid_Out & channel15_Kernel5_Valid_Out & channel16_Kernel5_Valid_Out & channel17_Kernel5_Valid_Out & channel18_Kernel5_Valid_Out & channel19_Kernel5_Valid_Out & channel20_Kernel5_Valid_Out & channel21_Kernel5_Valid_Out & channel22_Kernel5_Valid_Out & channel23_Kernel5_Valid_Out & channel24_Kernel5_Valid_Out & channel25_Kernel5_Valid_Out & channel26_Kernel5_Valid_Out & channel27_Kernel5_Valid_Out & channel28_Kernel5_Valid_Out & channel29_Kernel5_Valid_Out & channel30_Kernel5_Valid_Out & channel31_Kernel5_Valid_Out & channel32_Kernel5_Valid_Out & channel33_Kernel5_Valid_Out & channel34_Kernel5_Valid_Out & channel35_Kernel5_Valid_Out & channel36_Kernel5_Valid_Out & channel37_Kernel5_Valid_Out & channel38_Kernel5_Valid_Out & channel39_Kernel5_Valid_Out & channel40_Kernel5_Valid_Out & channel41_Kernel5_Valid_Out & channel42_Kernel5_Valid_Out & channel43_Kernel5_Valid_Out & channel44_Kernel5_Valid_Out & channel45_Kernel5_Valid_Out & channel46_Kernel5_Valid_Out & channel47_Kernel5_Valid_Out & channel48_Kernel5_Valid_Out & channel49_Kernel5_Valid_Out & channel50_Kernel5_Valid_Out & channel51_Kernel5_Valid_Out & channel52_Kernel5_Valid_Out & channel53_Kernel5_Valid_Out & channel54_Kernel5_Valid_Out & channel55_Kernel5_Valid_Out & channel56_Kernel5_Valid_Out & channel57_Kernel5_Valid_Out & channel58_Kernel5_Valid_Out & channel59_Kernel5_Valid_Out & channel60_Kernel5_Valid_Out & channel61_Kernel5_Valid_Out & channel62_Kernel5_Valid_Out & channel63_Kernel5_Valid_Out & channel64_Kernel5_Valid_Out;

	wire channel1_Kernel6_Valid_Out, channel2_Kernel6_Valid_Out, channel3_Kernel6_Valid_Out, channel4_Kernel6_Valid_Out, channel5_Kernel6_Valid_Out, channel6_Kernel6_Valid_Out, channel7_Kernel6_Valid_Out, channel8_Kernel6_Valid_Out, channel9_Kernel6_Valid_Out, channel10_Kernel6_Valid_Out, channel11_Kernel6_Valid_Out, channel12_Kernel6_Valid_Out, channel13_Kernel6_Valid_Out, channel14_Kernel6_Valid_Out, channel15_Kernel6_Valid_Out, channel16_Kernel6_Valid_Out, channel17_Kernel6_Valid_Out, channel18_Kernel6_Valid_Out, channel19_Kernel6_Valid_Out, channel20_Kernel6_Valid_Out, channel21_Kernel6_Valid_Out, channel22_Kernel6_Valid_Out, channel23_Kernel6_Valid_Out, channel24_Kernel6_Valid_Out, channel25_Kernel6_Valid_Out, channel26_Kernel6_Valid_Out, channel27_Kernel6_Valid_Out, channel28_Kernel6_Valid_Out, channel29_Kernel6_Valid_Out, channel30_Kernel6_Valid_Out, channel31_Kernel6_Valid_Out, channel32_Kernel6_Valid_Out, channel33_Kernel6_Valid_Out, channel34_Kernel6_Valid_Out, channel35_Kernel6_Valid_Out, channel36_Kernel6_Valid_Out, channel37_Kernel6_Valid_Out, channel38_Kernel6_Valid_Out, channel39_Kernel6_Valid_Out, channel40_Kernel6_Valid_Out, channel41_Kernel6_Valid_Out, channel42_Kernel6_Valid_Out, channel43_Kernel6_Valid_Out, channel44_Kernel6_Valid_Out, channel45_Kernel6_Valid_Out, channel46_Kernel6_Valid_Out, channel47_Kernel6_Valid_Out, channel48_Kernel6_Valid_Out, channel49_Kernel6_Valid_Out, channel50_Kernel6_Valid_Out, channel51_Kernel6_Valid_Out, channel52_Kernel6_Valid_Out, channel53_Kernel6_Valid_Out, channel54_Kernel6_Valid_Out, channel55_Kernel6_Valid_Out, channel56_Kernel6_Valid_Out, channel57_Kernel6_Valid_Out, channel58_Kernel6_Valid_Out, channel59_Kernel6_Valid_Out, channel60_Kernel6_Valid_Out, channel61_Kernel6_Valid_Out, channel62_Kernel6_Valid_Out, channel63_Kernel6_Valid_Out, channel64_Kernel6_Valid_Out;

	assign add_kernel6=channel1_Kernel6_Valid_Out & channel2_Kernel6_Valid_Out & channel3_Kernel6_Valid_Out & channel4_Kernel6_Valid_Out & channel5_Kernel6_Valid_Out & channel6_Kernel6_Valid_Out & channel7_Kernel6_Valid_Out & channel8_Kernel6_Valid_Out & channel9_Kernel6_Valid_Out & channel10_Kernel6_Valid_Out & channel11_Kernel6_Valid_Out & channel12_Kernel6_Valid_Out & channel13_Kernel6_Valid_Out & channel14_Kernel6_Valid_Out & channel15_Kernel6_Valid_Out & channel16_Kernel6_Valid_Out & channel17_Kernel6_Valid_Out & channel18_Kernel6_Valid_Out & channel19_Kernel6_Valid_Out & channel20_Kernel6_Valid_Out & channel21_Kernel6_Valid_Out & channel22_Kernel6_Valid_Out & channel23_Kernel6_Valid_Out & channel24_Kernel6_Valid_Out & channel25_Kernel6_Valid_Out & channel26_Kernel6_Valid_Out & channel27_Kernel6_Valid_Out & channel28_Kernel6_Valid_Out & channel29_Kernel6_Valid_Out & channel30_Kernel6_Valid_Out & channel31_Kernel6_Valid_Out & channel32_Kernel6_Valid_Out & channel33_Kernel6_Valid_Out & channel34_Kernel6_Valid_Out & channel35_Kernel6_Valid_Out & channel36_Kernel6_Valid_Out & channel37_Kernel6_Valid_Out & channel38_Kernel6_Valid_Out & channel39_Kernel6_Valid_Out & channel40_Kernel6_Valid_Out & channel41_Kernel6_Valid_Out & channel42_Kernel6_Valid_Out & channel43_Kernel6_Valid_Out & channel44_Kernel6_Valid_Out & channel45_Kernel6_Valid_Out & channel46_Kernel6_Valid_Out & channel47_Kernel6_Valid_Out & channel48_Kernel6_Valid_Out & channel49_Kernel6_Valid_Out & channel50_Kernel6_Valid_Out & channel51_Kernel6_Valid_Out & channel52_Kernel6_Valid_Out & channel53_Kernel6_Valid_Out & channel54_Kernel6_Valid_Out & channel55_Kernel6_Valid_Out & channel56_Kernel6_Valid_Out & channel57_Kernel6_Valid_Out & channel58_Kernel6_Valid_Out & channel59_Kernel6_Valid_Out & channel60_Kernel6_Valid_Out & channel61_Kernel6_Valid_Out & channel62_Kernel6_Valid_Out & channel63_Kernel6_Valid_Out & channel64_Kernel6_Valid_Out;

	wire channel1_Kernel7_Valid_Out, channel2_Kernel7_Valid_Out, channel3_Kernel7_Valid_Out, channel4_Kernel7_Valid_Out, channel5_Kernel7_Valid_Out, channel6_Kernel7_Valid_Out, channel7_Kernel7_Valid_Out, channel8_Kernel7_Valid_Out, channel9_Kernel7_Valid_Out, channel10_Kernel7_Valid_Out, channel11_Kernel7_Valid_Out, channel12_Kernel7_Valid_Out, channel13_Kernel7_Valid_Out, channel14_Kernel7_Valid_Out, channel15_Kernel7_Valid_Out, channel16_Kernel7_Valid_Out, channel17_Kernel7_Valid_Out, channel18_Kernel7_Valid_Out, channel19_Kernel7_Valid_Out, channel20_Kernel7_Valid_Out, channel21_Kernel7_Valid_Out, channel22_Kernel7_Valid_Out, channel23_Kernel7_Valid_Out, channel24_Kernel7_Valid_Out, channel25_Kernel7_Valid_Out, channel26_Kernel7_Valid_Out, channel27_Kernel7_Valid_Out, channel28_Kernel7_Valid_Out, channel29_Kernel7_Valid_Out, channel30_Kernel7_Valid_Out, channel31_Kernel7_Valid_Out, channel32_Kernel7_Valid_Out, channel33_Kernel7_Valid_Out, channel34_Kernel7_Valid_Out, channel35_Kernel7_Valid_Out, channel36_Kernel7_Valid_Out, channel37_Kernel7_Valid_Out, channel38_Kernel7_Valid_Out, channel39_Kernel7_Valid_Out, channel40_Kernel7_Valid_Out, channel41_Kernel7_Valid_Out, channel42_Kernel7_Valid_Out, channel43_Kernel7_Valid_Out, channel44_Kernel7_Valid_Out, channel45_Kernel7_Valid_Out, channel46_Kernel7_Valid_Out, channel47_Kernel7_Valid_Out, channel48_Kernel7_Valid_Out, channel49_Kernel7_Valid_Out, channel50_Kernel7_Valid_Out, channel51_Kernel7_Valid_Out, channel52_Kernel7_Valid_Out, channel53_Kernel7_Valid_Out, channel54_Kernel7_Valid_Out, channel55_Kernel7_Valid_Out, channel56_Kernel7_Valid_Out, channel57_Kernel7_Valid_Out, channel58_Kernel7_Valid_Out, channel59_Kernel7_Valid_Out, channel60_Kernel7_Valid_Out, channel61_Kernel7_Valid_Out, channel62_Kernel7_Valid_Out, channel63_Kernel7_Valid_Out, channel64_Kernel7_Valid_Out;

	assign add_kernel7=channel1_Kernel7_Valid_Out & channel2_Kernel7_Valid_Out & channel3_Kernel7_Valid_Out & channel4_Kernel7_Valid_Out & channel5_Kernel7_Valid_Out & channel6_Kernel7_Valid_Out & channel7_Kernel7_Valid_Out & channel8_Kernel7_Valid_Out & channel9_Kernel7_Valid_Out & channel10_Kernel7_Valid_Out & channel11_Kernel7_Valid_Out & channel12_Kernel7_Valid_Out & channel13_Kernel7_Valid_Out & channel14_Kernel7_Valid_Out & channel15_Kernel7_Valid_Out & channel16_Kernel7_Valid_Out & channel17_Kernel7_Valid_Out & channel18_Kernel7_Valid_Out & channel19_Kernel7_Valid_Out & channel20_Kernel7_Valid_Out & channel21_Kernel7_Valid_Out & channel22_Kernel7_Valid_Out & channel23_Kernel7_Valid_Out & channel24_Kernel7_Valid_Out & channel25_Kernel7_Valid_Out & channel26_Kernel7_Valid_Out & channel27_Kernel7_Valid_Out & channel28_Kernel7_Valid_Out & channel29_Kernel7_Valid_Out & channel30_Kernel7_Valid_Out & channel31_Kernel7_Valid_Out & channel32_Kernel7_Valid_Out & channel33_Kernel7_Valid_Out & channel34_Kernel7_Valid_Out & channel35_Kernel7_Valid_Out & channel36_Kernel7_Valid_Out & channel37_Kernel7_Valid_Out & channel38_Kernel7_Valid_Out & channel39_Kernel7_Valid_Out & channel40_Kernel7_Valid_Out & channel41_Kernel7_Valid_Out & channel42_Kernel7_Valid_Out & channel43_Kernel7_Valid_Out & channel44_Kernel7_Valid_Out & channel45_Kernel7_Valid_Out & channel46_Kernel7_Valid_Out & channel47_Kernel7_Valid_Out & channel48_Kernel7_Valid_Out & channel49_Kernel7_Valid_Out & channel50_Kernel7_Valid_Out & channel51_Kernel7_Valid_Out & channel52_Kernel7_Valid_Out & channel53_Kernel7_Valid_Out & channel54_Kernel7_Valid_Out & channel55_Kernel7_Valid_Out & channel56_Kernel7_Valid_Out & channel57_Kernel7_Valid_Out & channel58_Kernel7_Valid_Out & channel59_Kernel7_Valid_Out & channel60_Kernel7_Valid_Out & channel61_Kernel7_Valid_Out & channel62_Kernel7_Valid_Out & channel63_Kernel7_Valid_Out & channel64_Kernel7_Valid_Out;

	wire channel1_Kernel8_Valid_Out, channel2_Kernel8_Valid_Out, channel3_Kernel8_Valid_Out, channel4_Kernel8_Valid_Out, channel5_Kernel8_Valid_Out, channel6_Kernel8_Valid_Out, channel7_Kernel8_Valid_Out, channel8_Kernel8_Valid_Out, channel9_Kernel8_Valid_Out, channel10_Kernel8_Valid_Out, channel11_Kernel8_Valid_Out, channel12_Kernel8_Valid_Out, channel13_Kernel8_Valid_Out, channel14_Kernel8_Valid_Out, channel15_Kernel8_Valid_Out, channel16_Kernel8_Valid_Out, channel17_Kernel8_Valid_Out, channel18_Kernel8_Valid_Out, channel19_Kernel8_Valid_Out, channel20_Kernel8_Valid_Out, channel21_Kernel8_Valid_Out, channel22_Kernel8_Valid_Out, channel23_Kernel8_Valid_Out, channel24_Kernel8_Valid_Out, channel25_Kernel8_Valid_Out, channel26_Kernel8_Valid_Out, channel27_Kernel8_Valid_Out, channel28_Kernel8_Valid_Out, channel29_Kernel8_Valid_Out, channel30_Kernel8_Valid_Out, channel31_Kernel8_Valid_Out, channel32_Kernel8_Valid_Out, channel33_Kernel8_Valid_Out, channel34_Kernel8_Valid_Out, channel35_Kernel8_Valid_Out, channel36_Kernel8_Valid_Out, channel37_Kernel8_Valid_Out, channel38_Kernel8_Valid_Out, channel39_Kernel8_Valid_Out, channel40_Kernel8_Valid_Out, channel41_Kernel8_Valid_Out, channel42_Kernel8_Valid_Out, channel43_Kernel8_Valid_Out, channel44_Kernel8_Valid_Out, channel45_Kernel8_Valid_Out, channel46_Kernel8_Valid_Out, channel47_Kernel8_Valid_Out, channel48_Kernel8_Valid_Out, channel49_Kernel8_Valid_Out, channel50_Kernel8_Valid_Out, channel51_Kernel8_Valid_Out, channel52_Kernel8_Valid_Out, channel53_Kernel8_Valid_Out, channel54_Kernel8_Valid_Out, channel55_Kernel8_Valid_Out, channel56_Kernel8_Valid_Out, channel57_Kernel8_Valid_Out, channel58_Kernel8_Valid_Out, channel59_Kernel8_Valid_Out, channel60_Kernel8_Valid_Out, channel61_Kernel8_Valid_Out, channel62_Kernel8_Valid_Out, channel63_Kernel8_Valid_Out, channel64_Kernel8_Valid_Out;

	assign add_kernel8=channel1_Kernel8_Valid_Out & channel2_Kernel8_Valid_Out & channel3_Kernel8_Valid_Out & channel4_Kernel8_Valid_Out & channel5_Kernel8_Valid_Out & channel6_Kernel8_Valid_Out & channel7_Kernel8_Valid_Out & channel8_Kernel8_Valid_Out & channel9_Kernel8_Valid_Out & channel10_Kernel8_Valid_Out & channel11_Kernel8_Valid_Out & channel12_Kernel8_Valid_Out & channel13_Kernel8_Valid_Out & channel14_Kernel8_Valid_Out & channel15_Kernel8_Valid_Out & channel16_Kernel8_Valid_Out & channel17_Kernel8_Valid_Out & channel18_Kernel8_Valid_Out & channel19_Kernel8_Valid_Out & channel20_Kernel8_Valid_Out & channel21_Kernel8_Valid_Out & channel22_Kernel8_Valid_Out & channel23_Kernel8_Valid_Out & channel24_Kernel8_Valid_Out & channel25_Kernel8_Valid_Out & channel26_Kernel8_Valid_Out & channel27_Kernel8_Valid_Out & channel28_Kernel8_Valid_Out & channel29_Kernel8_Valid_Out & channel30_Kernel8_Valid_Out & channel31_Kernel8_Valid_Out & channel32_Kernel8_Valid_Out & channel33_Kernel8_Valid_Out & channel34_Kernel8_Valid_Out & channel35_Kernel8_Valid_Out & channel36_Kernel8_Valid_Out & channel37_Kernel8_Valid_Out & channel38_Kernel8_Valid_Out & channel39_Kernel8_Valid_Out & channel40_Kernel8_Valid_Out & channel41_Kernel8_Valid_Out & channel42_Kernel8_Valid_Out & channel43_Kernel8_Valid_Out & channel44_Kernel8_Valid_Out & channel45_Kernel8_Valid_Out & channel46_Kernel8_Valid_Out & channel47_Kernel8_Valid_Out & channel48_Kernel8_Valid_Out & channel49_Kernel8_Valid_Out & channel50_Kernel8_Valid_Out & channel51_Kernel8_Valid_Out & channel52_Kernel8_Valid_Out & channel53_Kernel8_Valid_Out & channel54_Kernel8_Valid_Out & channel55_Kernel8_Valid_Out & channel56_Kernel8_Valid_Out & channel57_Kernel8_Valid_Out & channel58_Kernel8_Valid_Out & channel59_Kernel8_Valid_Out & channel60_Kernel8_Valid_Out & channel61_Kernel8_Valid_Out & channel62_Kernel8_Valid_Out & channel63_Kernel8_Valid_Out & channel64_Kernel8_Valid_Out;

	wire channel1_Kernel9_Valid_Out, channel2_Kernel9_Valid_Out, channel3_Kernel9_Valid_Out, channel4_Kernel9_Valid_Out, channel5_Kernel9_Valid_Out, channel6_Kernel9_Valid_Out, channel7_Kernel9_Valid_Out, channel8_Kernel9_Valid_Out, channel9_Kernel9_Valid_Out, channel10_Kernel9_Valid_Out, channel11_Kernel9_Valid_Out, channel12_Kernel9_Valid_Out, channel13_Kernel9_Valid_Out, channel14_Kernel9_Valid_Out, channel15_Kernel9_Valid_Out, channel16_Kernel9_Valid_Out, channel17_Kernel9_Valid_Out, channel18_Kernel9_Valid_Out, channel19_Kernel9_Valid_Out, channel20_Kernel9_Valid_Out, channel21_Kernel9_Valid_Out, channel22_Kernel9_Valid_Out, channel23_Kernel9_Valid_Out, channel24_Kernel9_Valid_Out, channel25_Kernel9_Valid_Out, channel26_Kernel9_Valid_Out, channel27_Kernel9_Valid_Out, channel28_Kernel9_Valid_Out, channel29_Kernel9_Valid_Out, channel30_Kernel9_Valid_Out, channel31_Kernel9_Valid_Out, channel32_Kernel9_Valid_Out, channel33_Kernel9_Valid_Out, channel34_Kernel9_Valid_Out, channel35_Kernel9_Valid_Out, channel36_Kernel9_Valid_Out, channel37_Kernel9_Valid_Out, channel38_Kernel9_Valid_Out, channel39_Kernel9_Valid_Out, channel40_Kernel9_Valid_Out, channel41_Kernel9_Valid_Out, channel42_Kernel9_Valid_Out, channel43_Kernel9_Valid_Out, channel44_Kernel9_Valid_Out, channel45_Kernel9_Valid_Out, channel46_Kernel9_Valid_Out, channel47_Kernel9_Valid_Out, channel48_Kernel9_Valid_Out, channel49_Kernel9_Valid_Out, channel50_Kernel9_Valid_Out, channel51_Kernel9_Valid_Out, channel52_Kernel9_Valid_Out, channel53_Kernel9_Valid_Out, channel54_Kernel9_Valid_Out, channel55_Kernel9_Valid_Out, channel56_Kernel9_Valid_Out, channel57_Kernel9_Valid_Out, channel58_Kernel9_Valid_Out, channel59_Kernel9_Valid_Out, channel60_Kernel9_Valid_Out, channel61_Kernel9_Valid_Out, channel62_Kernel9_Valid_Out, channel63_Kernel9_Valid_Out, channel64_Kernel9_Valid_Out;

	assign add_kernel9=channel1_Kernel9_Valid_Out & channel2_Kernel9_Valid_Out & channel3_Kernel9_Valid_Out & channel4_Kernel9_Valid_Out & channel5_Kernel9_Valid_Out & channel6_Kernel9_Valid_Out & channel7_Kernel9_Valid_Out & channel8_Kernel9_Valid_Out & channel9_Kernel9_Valid_Out & channel10_Kernel9_Valid_Out & channel11_Kernel9_Valid_Out & channel12_Kernel9_Valid_Out & channel13_Kernel9_Valid_Out & channel14_Kernel9_Valid_Out & channel15_Kernel9_Valid_Out & channel16_Kernel9_Valid_Out & channel17_Kernel9_Valid_Out & channel18_Kernel9_Valid_Out & channel19_Kernel9_Valid_Out & channel20_Kernel9_Valid_Out & channel21_Kernel9_Valid_Out & channel22_Kernel9_Valid_Out & channel23_Kernel9_Valid_Out & channel24_Kernel9_Valid_Out & channel25_Kernel9_Valid_Out & channel26_Kernel9_Valid_Out & channel27_Kernel9_Valid_Out & channel28_Kernel9_Valid_Out & channel29_Kernel9_Valid_Out & channel30_Kernel9_Valid_Out & channel31_Kernel9_Valid_Out & channel32_Kernel9_Valid_Out & channel33_Kernel9_Valid_Out & channel34_Kernel9_Valid_Out & channel35_Kernel9_Valid_Out & channel36_Kernel9_Valid_Out & channel37_Kernel9_Valid_Out & channel38_Kernel9_Valid_Out & channel39_Kernel9_Valid_Out & channel40_Kernel9_Valid_Out & channel41_Kernel9_Valid_Out & channel42_Kernel9_Valid_Out & channel43_Kernel9_Valid_Out & channel44_Kernel9_Valid_Out & channel45_Kernel9_Valid_Out & channel46_Kernel9_Valid_Out & channel47_Kernel9_Valid_Out & channel48_Kernel9_Valid_Out & channel49_Kernel9_Valid_Out & channel50_Kernel9_Valid_Out & channel51_Kernel9_Valid_Out & channel52_Kernel9_Valid_Out & channel53_Kernel9_Valid_Out & channel54_Kernel9_Valid_Out & channel55_Kernel9_Valid_Out & channel56_Kernel9_Valid_Out & channel57_Kernel9_Valid_Out & channel58_Kernel9_Valid_Out & channel59_Kernel9_Valid_Out & channel60_Kernel9_Valid_Out & channel61_Kernel9_Valid_Out & channel62_Kernel9_Valid_Out & channel63_Kernel9_Valid_Out & channel64_Kernel9_Valid_Out;

	wire channel1_Kernel10_Valid_Out, channel2_Kernel10_Valid_Out, channel3_Kernel10_Valid_Out, channel4_Kernel10_Valid_Out, channel5_Kernel10_Valid_Out, channel6_Kernel10_Valid_Out, channel7_Kernel10_Valid_Out, channel8_Kernel10_Valid_Out, channel9_Kernel10_Valid_Out, channel10_Kernel10_Valid_Out, channel11_Kernel10_Valid_Out, channel12_Kernel10_Valid_Out, channel13_Kernel10_Valid_Out, channel14_Kernel10_Valid_Out, channel15_Kernel10_Valid_Out, channel16_Kernel10_Valid_Out, channel17_Kernel10_Valid_Out, channel18_Kernel10_Valid_Out, channel19_Kernel10_Valid_Out, channel20_Kernel10_Valid_Out, channel21_Kernel10_Valid_Out, channel22_Kernel10_Valid_Out, channel23_Kernel10_Valid_Out, channel24_Kernel10_Valid_Out, channel25_Kernel10_Valid_Out, channel26_Kernel10_Valid_Out, channel27_Kernel10_Valid_Out, channel28_Kernel10_Valid_Out, channel29_Kernel10_Valid_Out, channel30_Kernel10_Valid_Out, channel31_Kernel10_Valid_Out, channel32_Kernel10_Valid_Out, channel33_Kernel10_Valid_Out, channel34_Kernel10_Valid_Out, channel35_Kernel10_Valid_Out, channel36_Kernel10_Valid_Out, channel37_Kernel10_Valid_Out, channel38_Kernel10_Valid_Out, channel39_Kernel10_Valid_Out, channel40_Kernel10_Valid_Out, channel41_Kernel10_Valid_Out, channel42_Kernel10_Valid_Out, channel43_Kernel10_Valid_Out, channel44_Kernel10_Valid_Out, channel45_Kernel10_Valid_Out, channel46_Kernel10_Valid_Out, channel47_Kernel10_Valid_Out, channel48_Kernel10_Valid_Out, channel49_Kernel10_Valid_Out, channel50_Kernel10_Valid_Out, channel51_Kernel10_Valid_Out, channel52_Kernel10_Valid_Out, channel53_Kernel10_Valid_Out, channel54_Kernel10_Valid_Out, channel55_Kernel10_Valid_Out, channel56_Kernel10_Valid_Out, channel57_Kernel10_Valid_Out, channel58_Kernel10_Valid_Out, channel59_Kernel10_Valid_Out, channel60_Kernel10_Valid_Out, channel61_Kernel10_Valid_Out, channel62_Kernel10_Valid_Out, channel63_Kernel10_Valid_Out, channel64_Kernel10_Valid_Out;

	assign add_kernel10=channel1_Kernel10_Valid_Out & channel2_Kernel10_Valid_Out & channel3_Kernel10_Valid_Out & channel4_Kernel10_Valid_Out & channel5_Kernel10_Valid_Out & channel6_Kernel10_Valid_Out & channel7_Kernel10_Valid_Out & channel8_Kernel10_Valid_Out & channel9_Kernel10_Valid_Out & channel10_Kernel10_Valid_Out & channel11_Kernel10_Valid_Out & channel12_Kernel10_Valid_Out & channel13_Kernel10_Valid_Out & channel14_Kernel10_Valid_Out & channel15_Kernel10_Valid_Out & channel16_Kernel10_Valid_Out & channel17_Kernel10_Valid_Out & channel18_Kernel10_Valid_Out & channel19_Kernel10_Valid_Out & channel20_Kernel10_Valid_Out & channel21_Kernel10_Valid_Out & channel22_Kernel10_Valid_Out & channel23_Kernel10_Valid_Out & channel24_Kernel10_Valid_Out & channel25_Kernel10_Valid_Out & channel26_Kernel10_Valid_Out & channel27_Kernel10_Valid_Out & channel28_Kernel10_Valid_Out & channel29_Kernel10_Valid_Out & channel30_Kernel10_Valid_Out & channel31_Kernel10_Valid_Out & channel32_Kernel10_Valid_Out & channel33_Kernel10_Valid_Out & channel34_Kernel10_Valid_Out & channel35_Kernel10_Valid_Out & channel36_Kernel10_Valid_Out & channel37_Kernel10_Valid_Out & channel38_Kernel10_Valid_Out & channel39_Kernel10_Valid_Out & channel40_Kernel10_Valid_Out & channel41_Kernel10_Valid_Out & channel42_Kernel10_Valid_Out & channel43_Kernel10_Valid_Out & channel44_Kernel10_Valid_Out & channel45_Kernel10_Valid_Out & channel46_Kernel10_Valid_Out & channel47_Kernel10_Valid_Out & channel48_Kernel10_Valid_Out & channel49_Kernel10_Valid_Out & channel50_Kernel10_Valid_Out & channel51_Kernel10_Valid_Out & channel52_Kernel10_Valid_Out & channel53_Kernel10_Valid_Out & channel54_Kernel10_Valid_Out & channel55_Kernel10_Valid_Out & channel56_Kernel10_Valid_Out & channel57_Kernel10_Valid_Out & channel58_Kernel10_Valid_Out & channel59_Kernel10_Valid_Out & channel60_Kernel10_Valid_Out & channel61_Kernel10_Valid_Out & channel62_Kernel10_Valid_Out & channel63_Kernel10_Valid_Out & channel64_Kernel10_Valid_Out;

	wire channel1_Kernel11_Valid_Out, channel2_Kernel11_Valid_Out, channel3_Kernel11_Valid_Out, channel4_Kernel11_Valid_Out, channel5_Kernel11_Valid_Out, channel6_Kernel11_Valid_Out, channel7_Kernel11_Valid_Out, channel8_Kernel11_Valid_Out, channel9_Kernel11_Valid_Out, channel10_Kernel11_Valid_Out, channel11_Kernel11_Valid_Out, channel12_Kernel11_Valid_Out, channel13_Kernel11_Valid_Out, channel14_Kernel11_Valid_Out, channel15_Kernel11_Valid_Out, channel16_Kernel11_Valid_Out, channel17_Kernel11_Valid_Out, channel18_Kernel11_Valid_Out, channel19_Kernel11_Valid_Out, channel20_Kernel11_Valid_Out, channel21_Kernel11_Valid_Out, channel22_Kernel11_Valid_Out, channel23_Kernel11_Valid_Out, channel24_Kernel11_Valid_Out, channel25_Kernel11_Valid_Out, channel26_Kernel11_Valid_Out, channel27_Kernel11_Valid_Out, channel28_Kernel11_Valid_Out, channel29_Kernel11_Valid_Out, channel30_Kernel11_Valid_Out, channel31_Kernel11_Valid_Out, channel32_Kernel11_Valid_Out, channel33_Kernel11_Valid_Out, channel34_Kernel11_Valid_Out, channel35_Kernel11_Valid_Out, channel36_Kernel11_Valid_Out, channel37_Kernel11_Valid_Out, channel38_Kernel11_Valid_Out, channel39_Kernel11_Valid_Out, channel40_Kernel11_Valid_Out, channel41_Kernel11_Valid_Out, channel42_Kernel11_Valid_Out, channel43_Kernel11_Valid_Out, channel44_Kernel11_Valid_Out, channel45_Kernel11_Valid_Out, channel46_Kernel11_Valid_Out, channel47_Kernel11_Valid_Out, channel48_Kernel11_Valid_Out, channel49_Kernel11_Valid_Out, channel50_Kernel11_Valid_Out, channel51_Kernel11_Valid_Out, channel52_Kernel11_Valid_Out, channel53_Kernel11_Valid_Out, channel54_Kernel11_Valid_Out, channel55_Kernel11_Valid_Out, channel56_Kernel11_Valid_Out, channel57_Kernel11_Valid_Out, channel58_Kernel11_Valid_Out, channel59_Kernel11_Valid_Out, channel60_Kernel11_Valid_Out, channel61_Kernel11_Valid_Out, channel62_Kernel11_Valid_Out, channel63_Kernel11_Valid_Out, channel64_Kernel11_Valid_Out;

	assign add_kernel11=channel1_Kernel11_Valid_Out & channel2_Kernel11_Valid_Out & channel3_Kernel11_Valid_Out & channel4_Kernel11_Valid_Out & channel5_Kernel11_Valid_Out & channel6_Kernel11_Valid_Out & channel7_Kernel11_Valid_Out & channel8_Kernel11_Valid_Out & channel9_Kernel11_Valid_Out & channel10_Kernel11_Valid_Out & channel11_Kernel11_Valid_Out & channel12_Kernel11_Valid_Out & channel13_Kernel11_Valid_Out & channel14_Kernel11_Valid_Out & channel15_Kernel11_Valid_Out & channel16_Kernel11_Valid_Out & channel17_Kernel11_Valid_Out & channel18_Kernel11_Valid_Out & channel19_Kernel11_Valid_Out & channel20_Kernel11_Valid_Out & channel21_Kernel11_Valid_Out & channel22_Kernel11_Valid_Out & channel23_Kernel11_Valid_Out & channel24_Kernel11_Valid_Out & channel25_Kernel11_Valid_Out & channel26_Kernel11_Valid_Out & channel27_Kernel11_Valid_Out & channel28_Kernel11_Valid_Out & channel29_Kernel11_Valid_Out & channel30_Kernel11_Valid_Out & channel31_Kernel11_Valid_Out & channel32_Kernel11_Valid_Out & channel33_Kernel11_Valid_Out & channel34_Kernel11_Valid_Out & channel35_Kernel11_Valid_Out & channel36_Kernel11_Valid_Out & channel37_Kernel11_Valid_Out & channel38_Kernel11_Valid_Out & channel39_Kernel11_Valid_Out & channel40_Kernel11_Valid_Out & channel41_Kernel11_Valid_Out & channel42_Kernel11_Valid_Out & channel43_Kernel11_Valid_Out & channel44_Kernel11_Valid_Out & channel45_Kernel11_Valid_Out & channel46_Kernel11_Valid_Out & channel47_Kernel11_Valid_Out & channel48_Kernel11_Valid_Out & channel49_Kernel11_Valid_Out & channel50_Kernel11_Valid_Out & channel51_Kernel11_Valid_Out & channel52_Kernel11_Valid_Out & channel53_Kernel11_Valid_Out & channel54_Kernel11_Valid_Out & channel55_Kernel11_Valid_Out & channel56_Kernel11_Valid_Out & channel57_Kernel11_Valid_Out & channel58_Kernel11_Valid_Out & channel59_Kernel11_Valid_Out & channel60_Kernel11_Valid_Out & channel61_Kernel11_Valid_Out & channel62_Kernel11_Valid_Out & channel63_Kernel11_Valid_Out & channel64_Kernel11_Valid_Out;

	wire channel1_Kernel12_Valid_Out, channel2_Kernel12_Valid_Out, channel3_Kernel12_Valid_Out, channel4_Kernel12_Valid_Out, channel5_Kernel12_Valid_Out, channel6_Kernel12_Valid_Out, channel7_Kernel12_Valid_Out, channel8_Kernel12_Valid_Out, channel9_Kernel12_Valid_Out, channel10_Kernel12_Valid_Out, channel11_Kernel12_Valid_Out, channel12_Kernel12_Valid_Out, channel13_Kernel12_Valid_Out, channel14_Kernel12_Valid_Out, channel15_Kernel12_Valid_Out, channel16_Kernel12_Valid_Out, channel17_Kernel12_Valid_Out, channel18_Kernel12_Valid_Out, channel19_Kernel12_Valid_Out, channel20_Kernel12_Valid_Out, channel21_Kernel12_Valid_Out, channel22_Kernel12_Valid_Out, channel23_Kernel12_Valid_Out, channel24_Kernel12_Valid_Out, channel25_Kernel12_Valid_Out, channel26_Kernel12_Valid_Out, channel27_Kernel12_Valid_Out, channel28_Kernel12_Valid_Out, channel29_Kernel12_Valid_Out, channel30_Kernel12_Valid_Out, channel31_Kernel12_Valid_Out, channel32_Kernel12_Valid_Out, channel33_Kernel12_Valid_Out, channel34_Kernel12_Valid_Out, channel35_Kernel12_Valid_Out, channel36_Kernel12_Valid_Out, channel37_Kernel12_Valid_Out, channel38_Kernel12_Valid_Out, channel39_Kernel12_Valid_Out, channel40_Kernel12_Valid_Out, channel41_Kernel12_Valid_Out, channel42_Kernel12_Valid_Out, channel43_Kernel12_Valid_Out, channel44_Kernel12_Valid_Out, channel45_Kernel12_Valid_Out, channel46_Kernel12_Valid_Out, channel47_Kernel12_Valid_Out, channel48_Kernel12_Valid_Out, channel49_Kernel12_Valid_Out, channel50_Kernel12_Valid_Out, channel51_Kernel12_Valid_Out, channel52_Kernel12_Valid_Out, channel53_Kernel12_Valid_Out, channel54_Kernel12_Valid_Out, channel55_Kernel12_Valid_Out, channel56_Kernel12_Valid_Out, channel57_Kernel12_Valid_Out, channel58_Kernel12_Valid_Out, channel59_Kernel12_Valid_Out, channel60_Kernel12_Valid_Out, channel61_Kernel12_Valid_Out, channel62_Kernel12_Valid_Out, channel63_Kernel12_Valid_Out, channel64_Kernel12_Valid_Out;

	assign add_kernel12=channel1_Kernel12_Valid_Out & channel2_Kernel12_Valid_Out & channel3_Kernel12_Valid_Out & channel4_Kernel12_Valid_Out & channel5_Kernel12_Valid_Out & channel6_Kernel12_Valid_Out & channel7_Kernel12_Valid_Out & channel8_Kernel12_Valid_Out & channel9_Kernel12_Valid_Out & channel10_Kernel12_Valid_Out & channel11_Kernel12_Valid_Out & channel12_Kernel12_Valid_Out & channel13_Kernel12_Valid_Out & channel14_Kernel12_Valid_Out & channel15_Kernel12_Valid_Out & channel16_Kernel12_Valid_Out & channel17_Kernel12_Valid_Out & channel18_Kernel12_Valid_Out & channel19_Kernel12_Valid_Out & channel20_Kernel12_Valid_Out & channel21_Kernel12_Valid_Out & channel22_Kernel12_Valid_Out & channel23_Kernel12_Valid_Out & channel24_Kernel12_Valid_Out & channel25_Kernel12_Valid_Out & channel26_Kernel12_Valid_Out & channel27_Kernel12_Valid_Out & channel28_Kernel12_Valid_Out & channel29_Kernel12_Valid_Out & channel30_Kernel12_Valid_Out & channel31_Kernel12_Valid_Out & channel32_Kernel12_Valid_Out & channel33_Kernel12_Valid_Out & channel34_Kernel12_Valid_Out & channel35_Kernel12_Valid_Out & channel36_Kernel12_Valid_Out & channel37_Kernel12_Valid_Out & channel38_Kernel12_Valid_Out & channel39_Kernel12_Valid_Out & channel40_Kernel12_Valid_Out & channel41_Kernel12_Valid_Out & channel42_Kernel12_Valid_Out & channel43_Kernel12_Valid_Out & channel44_Kernel12_Valid_Out & channel45_Kernel12_Valid_Out & channel46_Kernel12_Valid_Out & channel47_Kernel12_Valid_Out & channel48_Kernel12_Valid_Out & channel49_Kernel12_Valid_Out & channel50_Kernel12_Valid_Out & channel51_Kernel12_Valid_Out & channel52_Kernel12_Valid_Out & channel53_Kernel12_Valid_Out & channel54_Kernel12_Valid_Out & channel55_Kernel12_Valid_Out & channel56_Kernel12_Valid_Out & channel57_Kernel12_Valid_Out & channel58_Kernel12_Valid_Out & channel59_Kernel12_Valid_Out & channel60_Kernel12_Valid_Out & channel61_Kernel12_Valid_Out & channel62_Kernel12_Valid_Out & channel63_Kernel12_Valid_Out & channel64_Kernel12_Valid_Out;

	wire channel1_Kernel13_Valid_Out, channel2_Kernel13_Valid_Out, channel3_Kernel13_Valid_Out, channel4_Kernel13_Valid_Out, channel5_Kernel13_Valid_Out, channel6_Kernel13_Valid_Out, channel7_Kernel13_Valid_Out, channel8_Kernel13_Valid_Out, channel9_Kernel13_Valid_Out, channel10_Kernel13_Valid_Out, channel11_Kernel13_Valid_Out, channel12_Kernel13_Valid_Out, channel13_Kernel13_Valid_Out, channel14_Kernel13_Valid_Out, channel15_Kernel13_Valid_Out, channel16_Kernel13_Valid_Out, channel17_Kernel13_Valid_Out, channel18_Kernel13_Valid_Out, channel19_Kernel13_Valid_Out, channel20_Kernel13_Valid_Out, channel21_Kernel13_Valid_Out, channel22_Kernel13_Valid_Out, channel23_Kernel13_Valid_Out, channel24_Kernel13_Valid_Out, channel25_Kernel13_Valid_Out, channel26_Kernel13_Valid_Out, channel27_Kernel13_Valid_Out, channel28_Kernel13_Valid_Out, channel29_Kernel13_Valid_Out, channel30_Kernel13_Valid_Out, channel31_Kernel13_Valid_Out, channel32_Kernel13_Valid_Out, channel33_Kernel13_Valid_Out, channel34_Kernel13_Valid_Out, channel35_Kernel13_Valid_Out, channel36_Kernel13_Valid_Out, channel37_Kernel13_Valid_Out, channel38_Kernel13_Valid_Out, channel39_Kernel13_Valid_Out, channel40_Kernel13_Valid_Out, channel41_Kernel13_Valid_Out, channel42_Kernel13_Valid_Out, channel43_Kernel13_Valid_Out, channel44_Kernel13_Valid_Out, channel45_Kernel13_Valid_Out, channel46_Kernel13_Valid_Out, channel47_Kernel13_Valid_Out, channel48_Kernel13_Valid_Out, channel49_Kernel13_Valid_Out, channel50_Kernel13_Valid_Out, channel51_Kernel13_Valid_Out, channel52_Kernel13_Valid_Out, channel53_Kernel13_Valid_Out, channel54_Kernel13_Valid_Out, channel55_Kernel13_Valid_Out, channel56_Kernel13_Valid_Out, channel57_Kernel13_Valid_Out, channel58_Kernel13_Valid_Out, channel59_Kernel13_Valid_Out, channel60_Kernel13_Valid_Out, channel61_Kernel13_Valid_Out, channel62_Kernel13_Valid_Out, channel63_Kernel13_Valid_Out, channel64_Kernel13_Valid_Out;

	assign add_kernel13=channel1_Kernel13_Valid_Out & channel2_Kernel13_Valid_Out & channel3_Kernel13_Valid_Out & channel4_Kernel13_Valid_Out & channel5_Kernel13_Valid_Out & channel6_Kernel13_Valid_Out & channel7_Kernel13_Valid_Out & channel8_Kernel13_Valid_Out & channel9_Kernel13_Valid_Out & channel10_Kernel13_Valid_Out & channel11_Kernel13_Valid_Out & channel12_Kernel13_Valid_Out & channel13_Kernel13_Valid_Out & channel14_Kernel13_Valid_Out & channel15_Kernel13_Valid_Out & channel16_Kernel13_Valid_Out & channel17_Kernel13_Valid_Out & channel18_Kernel13_Valid_Out & channel19_Kernel13_Valid_Out & channel20_Kernel13_Valid_Out & channel21_Kernel13_Valid_Out & channel22_Kernel13_Valid_Out & channel23_Kernel13_Valid_Out & channel24_Kernel13_Valid_Out & channel25_Kernel13_Valid_Out & channel26_Kernel13_Valid_Out & channel27_Kernel13_Valid_Out & channel28_Kernel13_Valid_Out & channel29_Kernel13_Valid_Out & channel30_Kernel13_Valid_Out & channel31_Kernel13_Valid_Out & channel32_Kernel13_Valid_Out & channel33_Kernel13_Valid_Out & channel34_Kernel13_Valid_Out & channel35_Kernel13_Valid_Out & channel36_Kernel13_Valid_Out & channel37_Kernel13_Valid_Out & channel38_Kernel13_Valid_Out & channel39_Kernel13_Valid_Out & channel40_Kernel13_Valid_Out & channel41_Kernel13_Valid_Out & channel42_Kernel13_Valid_Out & channel43_Kernel13_Valid_Out & channel44_Kernel13_Valid_Out & channel45_Kernel13_Valid_Out & channel46_Kernel13_Valid_Out & channel47_Kernel13_Valid_Out & channel48_Kernel13_Valid_Out & channel49_Kernel13_Valid_Out & channel50_Kernel13_Valid_Out & channel51_Kernel13_Valid_Out & channel52_Kernel13_Valid_Out & channel53_Kernel13_Valid_Out & channel54_Kernel13_Valid_Out & channel55_Kernel13_Valid_Out & channel56_Kernel13_Valid_Out & channel57_Kernel13_Valid_Out & channel58_Kernel13_Valid_Out & channel59_Kernel13_Valid_Out & channel60_Kernel13_Valid_Out & channel61_Kernel13_Valid_Out & channel62_Kernel13_Valid_Out & channel63_Kernel13_Valid_Out & channel64_Kernel13_Valid_Out;

	wire channel1_Kernel14_Valid_Out, channel2_Kernel14_Valid_Out, channel3_Kernel14_Valid_Out, channel4_Kernel14_Valid_Out, channel5_Kernel14_Valid_Out, channel6_Kernel14_Valid_Out, channel7_Kernel14_Valid_Out, channel8_Kernel14_Valid_Out, channel9_Kernel14_Valid_Out, channel10_Kernel14_Valid_Out, channel11_Kernel14_Valid_Out, channel12_Kernel14_Valid_Out, channel13_Kernel14_Valid_Out, channel14_Kernel14_Valid_Out, channel15_Kernel14_Valid_Out, channel16_Kernel14_Valid_Out, channel17_Kernel14_Valid_Out, channel18_Kernel14_Valid_Out, channel19_Kernel14_Valid_Out, channel20_Kernel14_Valid_Out, channel21_Kernel14_Valid_Out, channel22_Kernel14_Valid_Out, channel23_Kernel14_Valid_Out, channel24_Kernel14_Valid_Out, channel25_Kernel14_Valid_Out, channel26_Kernel14_Valid_Out, channel27_Kernel14_Valid_Out, channel28_Kernel14_Valid_Out, channel29_Kernel14_Valid_Out, channel30_Kernel14_Valid_Out, channel31_Kernel14_Valid_Out, channel32_Kernel14_Valid_Out, channel33_Kernel14_Valid_Out, channel34_Kernel14_Valid_Out, channel35_Kernel14_Valid_Out, channel36_Kernel14_Valid_Out, channel37_Kernel14_Valid_Out, channel38_Kernel14_Valid_Out, channel39_Kernel14_Valid_Out, channel40_Kernel14_Valid_Out, channel41_Kernel14_Valid_Out, channel42_Kernel14_Valid_Out, channel43_Kernel14_Valid_Out, channel44_Kernel14_Valid_Out, channel45_Kernel14_Valid_Out, channel46_Kernel14_Valid_Out, channel47_Kernel14_Valid_Out, channel48_Kernel14_Valid_Out, channel49_Kernel14_Valid_Out, channel50_Kernel14_Valid_Out, channel51_Kernel14_Valid_Out, channel52_Kernel14_Valid_Out, channel53_Kernel14_Valid_Out, channel54_Kernel14_Valid_Out, channel55_Kernel14_Valid_Out, channel56_Kernel14_Valid_Out, channel57_Kernel14_Valid_Out, channel58_Kernel14_Valid_Out, channel59_Kernel14_Valid_Out, channel60_Kernel14_Valid_Out, channel61_Kernel14_Valid_Out, channel62_Kernel14_Valid_Out, channel63_Kernel14_Valid_Out, channel64_Kernel14_Valid_Out;

	assign add_kernel14=channel1_Kernel14_Valid_Out & channel2_Kernel14_Valid_Out & channel3_Kernel14_Valid_Out & channel4_Kernel14_Valid_Out & channel5_Kernel14_Valid_Out & channel6_Kernel14_Valid_Out & channel7_Kernel14_Valid_Out & channel8_Kernel14_Valid_Out & channel9_Kernel14_Valid_Out & channel10_Kernel14_Valid_Out & channel11_Kernel14_Valid_Out & channel12_Kernel14_Valid_Out & channel13_Kernel14_Valid_Out & channel14_Kernel14_Valid_Out & channel15_Kernel14_Valid_Out & channel16_Kernel14_Valid_Out & channel17_Kernel14_Valid_Out & channel18_Kernel14_Valid_Out & channel19_Kernel14_Valid_Out & channel20_Kernel14_Valid_Out & channel21_Kernel14_Valid_Out & channel22_Kernel14_Valid_Out & channel23_Kernel14_Valid_Out & channel24_Kernel14_Valid_Out & channel25_Kernel14_Valid_Out & channel26_Kernel14_Valid_Out & channel27_Kernel14_Valid_Out & channel28_Kernel14_Valid_Out & channel29_Kernel14_Valid_Out & channel30_Kernel14_Valid_Out & channel31_Kernel14_Valid_Out & channel32_Kernel14_Valid_Out & channel33_Kernel14_Valid_Out & channel34_Kernel14_Valid_Out & channel35_Kernel14_Valid_Out & channel36_Kernel14_Valid_Out & channel37_Kernel14_Valid_Out & channel38_Kernel14_Valid_Out & channel39_Kernel14_Valid_Out & channel40_Kernel14_Valid_Out & channel41_Kernel14_Valid_Out & channel42_Kernel14_Valid_Out & channel43_Kernel14_Valid_Out & channel44_Kernel14_Valid_Out & channel45_Kernel14_Valid_Out & channel46_Kernel14_Valid_Out & channel47_Kernel14_Valid_Out & channel48_Kernel14_Valid_Out & channel49_Kernel14_Valid_Out & channel50_Kernel14_Valid_Out & channel51_Kernel14_Valid_Out & channel52_Kernel14_Valid_Out & channel53_Kernel14_Valid_Out & channel54_Kernel14_Valid_Out & channel55_Kernel14_Valid_Out & channel56_Kernel14_Valid_Out & channel57_Kernel14_Valid_Out & channel58_Kernel14_Valid_Out & channel59_Kernel14_Valid_Out & channel60_Kernel14_Valid_Out & channel61_Kernel14_Valid_Out & channel62_Kernel14_Valid_Out & channel63_Kernel14_Valid_Out & channel64_Kernel14_Valid_Out;

	wire channel1_Kernel15_Valid_Out, channel2_Kernel15_Valid_Out, channel3_Kernel15_Valid_Out, channel4_Kernel15_Valid_Out, channel5_Kernel15_Valid_Out, channel6_Kernel15_Valid_Out, channel7_Kernel15_Valid_Out, channel8_Kernel15_Valid_Out, channel9_Kernel15_Valid_Out, channel10_Kernel15_Valid_Out, channel11_Kernel15_Valid_Out, channel12_Kernel15_Valid_Out, channel13_Kernel15_Valid_Out, channel14_Kernel15_Valid_Out, channel15_Kernel15_Valid_Out, channel16_Kernel15_Valid_Out, channel17_Kernel15_Valid_Out, channel18_Kernel15_Valid_Out, channel19_Kernel15_Valid_Out, channel20_Kernel15_Valid_Out, channel21_Kernel15_Valid_Out, channel22_Kernel15_Valid_Out, channel23_Kernel15_Valid_Out, channel24_Kernel15_Valid_Out, channel25_Kernel15_Valid_Out, channel26_Kernel15_Valid_Out, channel27_Kernel15_Valid_Out, channel28_Kernel15_Valid_Out, channel29_Kernel15_Valid_Out, channel30_Kernel15_Valid_Out, channel31_Kernel15_Valid_Out, channel32_Kernel15_Valid_Out, channel33_Kernel15_Valid_Out, channel34_Kernel15_Valid_Out, channel35_Kernel15_Valid_Out, channel36_Kernel15_Valid_Out, channel37_Kernel15_Valid_Out, channel38_Kernel15_Valid_Out, channel39_Kernel15_Valid_Out, channel40_Kernel15_Valid_Out, channel41_Kernel15_Valid_Out, channel42_Kernel15_Valid_Out, channel43_Kernel15_Valid_Out, channel44_Kernel15_Valid_Out, channel45_Kernel15_Valid_Out, channel46_Kernel15_Valid_Out, channel47_Kernel15_Valid_Out, channel48_Kernel15_Valid_Out, channel49_Kernel15_Valid_Out, channel50_Kernel15_Valid_Out, channel51_Kernel15_Valid_Out, channel52_Kernel15_Valid_Out, channel53_Kernel15_Valid_Out, channel54_Kernel15_Valid_Out, channel55_Kernel15_Valid_Out, channel56_Kernel15_Valid_Out, channel57_Kernel15_Valid_Out, channel58_Kernel15_Valid_Out, channel59_Kernel15_Valid_Out, channel60_Kernel15_Valid_Out, channel61_Kernel15_Valid_Out, channel62_Kernel15_Valid_Out, channel63_Kernel15_Valid_Out, channel64_Kernel15_Valid_Out;

	assign add_kernel15=channel1_Kernel15_Valid_Out & channel2_Kernel15_Valid_Out & channel3_Kernel15_Valid_Out & channel4_Kernel15_Valid_Out & channel5_Kernel15_Valid_Out & channel6_Kernel15_Valid_Out & channel7_Kernel15_Valid_Out & channel8_Kernel15_Valid_Out & channel9_Kernel15_Valid_Out & channel10_Kernel15_Valid_Out & channel11_Kernel15_Valid_Out & channel12_Kernel15_Valid_Out & channel13_Kernel15_Valid_Out & channel14_Kernel15_Valid_Out & channel15_Kernel15_Valid_Out & channel16_Kernel15_Valid_Out & channel17_Kernel15_Valid_Out & channel18_Kernel15_Valid_Out & channel19_Kernel15_Valid_Out & channel20_Kernel15_Valid_Out & channel21_Kernel15_Valid_Out & channel22_Kernel15_Valid_Out & channel23_Kernel15_Valid_Out & channel24_Kernel15_Valid_Out & channel25_Kernel15_Valid_Out & channel26_Kernel15_Valid_Out & channel27_Kernel15_Valid_Out & channel28_Kernel15_Valid_Out & channel29_Kernel15_Valid_Out & channel30_Kernel15_Valid_Out & channel31_Kernel15_Valid_Out & channel32_Kernel15_Valid_Out & channel33_Kernel15_Valid_Out & channel34_Kernel15_Valid_Out & channel35_Kernel15_Valid_Out & channel36_Kernel15_Valid_Out & channel37_Kernel15_Valid_Out & channel38_Kernel15_Valid_Out & channel39_Kernel15_Valid_Out & channel40_Kernel15_Valid_Out & channel41_Kernel15_Valid_Out & channel42_Kernel15_Valid_Out & channel43_Kernel15_Valid_Out & channel44_Kernel15_Valid_Out & channel45_Kernel15_Valid_Out & channel46_Kernel15_Valid_Out & channel47_Kernel15_Valid_Out & channel48_Kernel15_Valid_Out & channel49_Kernel15_Valid_Out & channel50_Kernel15_Valid_Out & channel51_Kernel15_Valid_Out & channel52_Kernel15_Valid_Out & channel53_Kernel15_Valid_Out & channel54_Kernel15_Valid_Out & channel55_Kernel15_Valid_Out & channel56_Kernel15_Valid_Out & channel57_Kernel15_Valid_Out & channel58_Kernel15_Valid_Out & channel59_Kernel15_Valid_Out & channel60_Kernel15_Valid_Out & channel61_Kernel15_Valid_Out & channel62_Kernel15_Valid_Out & channel63_Kernel15_Valid_Out & channel64_Kernel15_Valid_Out;

	wire channel1_Kernel16_Valid_Out, channel2_Kernel16_Valid_Out, channel3_Kernel16_Valid_Out, channel4_Kernel16_Valid_Out, channel5_Kernel16_Valid_Out, channel6_Kernel16_Valid_Out, channel7_Kernel16_Valid_Out, channel8_Kernel16_Valid_Out, channel9_Kernel16_Valid_Out, channel10_Kernel16_Valid_Out, channel11_Kernel16_Valid_Out, channel12_Kernel16_Valid_Out, channel13_Kernel16_Valid_Out, channel14_Kernel16_Valid_Out, channel15_Kernel16_Valid_Out, channel16_Kernel16_Valid_Out, channel17_Kernel16_Valid_Out, channel18_Kernel16_Valid_Out, channel19_Kernel16_Valid_Out, channel20_Kernel16_Valid_Out, channel21_Kernel16_Valid_Out, channel22_Kernel16_Valid_Out, channel23_Kernel16_Valid_Out, channel24_Kernel16_Valid_Out, channel25_Kernel16_Valid_Out, channel26_Kernel16_Valid_Out, channel27_Kernel16_Valid_Out, channel28_Kernel16_Valid_Out, channel29_Kernel16_Valid_Out, channel30_Kernel16_Valid_Out, channel31_Kernel16_Valid_Out, channel32_Kernel16_Valid_Out, channel33_Kernel16_Valid_Out, channel34_Kernel16_Valid_Out, channel35_Kernel16_Valid_Out, channel36_Kernel16_Valid_Out, channel37_Kernel16_Valid_Out, channel38_Kernel16_Valid_Out, channel39_Kernel16_Valid_Out, channel40_Kernel16_Valid_Out, channel41_Kernel16_Valid_Out, channel42_Kernel16_Valid_Out, channel43_Kernel16_Valid_Out, channel44_Kernel16_Valid_Out, channel45_Kernel16_Valid_Out, channel46_Kernel16_Valid_Out, channel47_Kernel16_Valid_Out, channel48_Kernel16_Valid_Out, channel49_Kernel16_Valid_Out, channel50_Kernel16_Valid_Out, channel51_Kernel16_Valid_Out, channel52_Kernel16_Valid_Out, channel53_Kernel16_Valid_Out, channel54_Kernel16_Valid_Out, channel55_Kernel16_Valid_Out, channel56_Kernel16_Valid_Out, channel57_Kernel16_Valid_Out, channel58_Kernel16_Valid_Out, channel59_Kernel16_Valid_Out, channel60_Kernel16_Valid_Out, channel61_Kernel16_Valid_Out, channel62_Kernel16_Valid_Out, channel63_Kernel16_Valid_Out, channel64_Kernel16_Valid_Out;

	assign add_kernel16=channel1_Kernel16_Valid_Out & channel2_Kernel16_Valid_Out & channel3_Kernel16_Valid_Out & channel4_Kernel16_Valid_Out & channel5_Kernel16_Valid_Out & channel6_Kernel16_Valid_Out & channel7_Kernel16_Valid_Out & channel8_Kernel16_Valid_Out & channel9_Kernel16_Valid_Out & channel10_Kernel16_Valid_Out & channel11_Kernel16_Valid_Out & channel12_Kernel16_Valid_Out & channel13_Kernel16_Valid_Out & channel14_Kernel16_Valid_Out & channel15_Kernel16_Valid_Out & channel16_Kernel16_Valid_Out & channel17_Kernel16_Valid_Out & channel18_Kernel16_Valid_Out & channel19_Kernel16_Valid_Out & channel20_Kernel16_Valid_Out & channel21_Kernel16_Valid_Out & channel22_Kernel16_Valid_Out & channel23_Kernel16_Valid_Out & channel24_Kernel16_Valid_Out & channel25_Kernel16_Valid_Out & channel26_Kernel16_Valid_Out & channel27_Kernel16_Valid_Out & channel28_Kernel16_Valid_Out & channel29_Kernel16_Valid_Out & channel30_Kernel16_Valid_Out & channel31_Kernel16_Valid_Out & channel32_Kernel16_Valid_Out & channel33_Kernel16_Valid_Out & channel34_Kernel16_Valid_Out & channel35_Kernel16_Valid_Out & channel36_Kernel16_Valid_Out & channel37_Kernel16_Valid_Out & channel38_Kernel16_Valid_Out & channel39_Kernel16_Valid_Out & channel40_Kernel16_Valid_Out & channel41_Kernel16_Valid_Out & channel42_Kernel16_Valid_Out & channel43_Kernel16_Valid_Out & channel44_Kernel16_Valid_Out & channel45_Kernel16_Valid_Out & channel46_Kernel16_Valid_Out & channel47_Kernel16_Valid_Out & channel48_Kernel16_Valid_Out & channel49_Kernel16_Valid_Out & channel50_Kernel16_Valid_Out & channel51_Kernel16_Valid_Out & channel52_Kernel16_Valid_Out & channel53_Kernel16_Valid_Out & channel54_Kernel16_Valid_Out & channel55_Kernel16_Valid_Out & channel56_Kernel16_Valid_Out & channel57_Kernel16_Valid_Out & channel58_Kernel16_Valid_Out & channel59_Kernel16_Valid_Out & channel60_Kernel16_Valid_Out & channel61_Kernel16_Valid_Out & channel62_Kernel16_Valid_Out & channel63_Kernel16_Valid_Out & channel64_Kernel16_Valid_Out;

	wire channel1_Kernel17_Valid_Out, channel2_Kernel17_Valid_Out, channel3_Kernel17_Valid_Out, channel4_Kernel17_Valid_Out, channel5_Kernel17_Valid_Out, channel6_Kernel17_Valid_Out, channel7_Kernel17_Valid_Out, channel8_Kernel17_Valid_Out, channel9_Kernel17_Valid_Out, channel10_Kernel17_Valid_Out, channel11_Kernel17_Valid_Out, channel12_Kernel17_Valid_Out, channel13_Kernel17_Valid_Out, channel14_Kernel17_Valid_Out, channel15_Kernel17_Valid_Out, channel16_Kernel17_Valid_Out, channel17_Kernel17_Valid_Out, channel18_Kernel17_Valid_Out, channel19_Kernel17_Valid_Out, channel20_Kernel17_Valid_Out, channel21_Kernel17_Valid_Out, channel22_Kernel17_Valid_Out, channel23_Kernel17_Valid_Out, channel24_Kernel17_Valid_Out, channel25_Kernel17_Valid_Out, channel26_Kernel17_Valid_Out, channel27_Kernel17_Valid_Out, channel28_Kernel17_Valid_Out, channel29_Kernel17_Valid_Out, channel30_Kernel17_Valid_Out, channel31_Kernel17_Valid_Out, channel32_Kernel17_Valid_Out, channel33_Kernel17_Valid_Out, channel34_Kernel17_Valid_Out, channel35_Kernel17_Valid_Out, channel36_Kernel17_Valid_Out, channel37_Kernel17_Valid_Out, channel38_Kernel17_Valid_Out, channel39_Kernel17_Valid_Out, channel40_Kernel17_Valid_Out, channel41_Kernel17_Valid_Out, channel42_Kernel17_Valid_Out, channel43_Kernel17_Valid_Out, channel44_Kernel17_Valid_Out, channel45_Kernel17_Valid_Out, channel46_Kernel17_Valid_Out, channel47_Kernel17_Valid_Out, channel48_Kernel17_Valid_Out, channel49_Kernel17_Valid_Out, channel50_Kernel17_Valid_Out, channel51_Kernel17_Valid_Out, channel52_Kernel17_Valid_Out, channel53_Kernel17_Valid_Out, channel54_Kernel17_Valid_Out, channel55_Kernel17_Valid_Out, channel56_Kernel17_Valid_Out, channel57_Kernel17_Valid_Out, channel58_Kernel17_Valid_Out, channel59_Kernel17_Valid_Out, channel60_Kernel17_Valid_Out, channel61_Kernel17_Valid_Out, channel62_Kernel17_Valid_Out, channel63_Kernel17_Valid_Out, channel64_Kernel17_Valid_Out;

	assign add_kernel17=channel1_Kernel17_Valid_Out & channel2_Kernel17_Valid_Out & channel3_Kernel17_Valid_Out & channel4_Kernel17_Valid_Out & channel5_Kernel17_Valid_Out & channel6_Kernel17_Valid_Out & channel7_Kernel17_Valid_Out & channel8_Kernel17_Valid_Out & channel9_Kernel17_Valid_Out & channel10_Kernel17_Valid_Out & channel11_Kernel17_Valid_Out & channel12_Kernel17_Valid_Out & channel13_Kernel17_Valid_Out & channel14_Kernel17_Valid_Out & channel15_Kernel17_Valid_Out & channel16_Kernel17_Valid_Out & channel17_Kernel17_Valid_Out & channel18_Kernel17_Valid_Out & channel19_Kernel17_Valid_Out & channel20_Kernel17_Valid_Out & channel21_Kernel17_Valid_Out & channel22_Kernel17_Valid_Out & channel23_Kernel17_Valid_Out & channel24_Kernel17_Valid_Out & channel25_Kernel17_Valid_Out & channel26_Kernel17_Valid_Out & channel27_Kernel17_Valid_Out & channel28_Kernel17_Valid_Out & channel29_Kernel17_Valid_Out & channel30_Kernel17_Valid_Out & channel31_Kernel17_Valid_Out & channel32_Kernel17_Valid_Out & channel33_Kernel17_Valid_Out & channel34_Kernel17_Valid_Out & channel35_Kernel17_Valid_Out & channel36_Kernel17_Valid_Out & channel37_Kernel17_Valid_Out & channel38_Kernel17_Valid_Out & channel39_Kernel17_Valid_Out & channel40_Kernel17_Valid_Out & channel41_Kernel17_Valid_Out & channel42_Kernel17_Valid_Out & channel43_Kernel17_Valid_Out & channel44_Kernel17_Valid_Out & channel45_Kernel17_Valid_Out & channel46_Kernel17_Valid_Out & channel47_Kernel17_Valid_Out & channel48_Kernel17_Valid_Out & channel49_Kernel17_Valid_Out & channel50_Kernel17_Valid_Out & channel51_Kernel17_Valid_Out & channel52_Kernel17_Valid_Out & channel53_Kernel17_Valid_Out & channel54_Kernel17_Valid_Out & channel55_Kernel17_Valid_Out & channel56_Kernel17_Valid_Out & channel57_Kernel17_Valid_Out & channel58_Kernel17_Valid_Out & channel59_Kernel17_Valid_Out & channel60_Kernel17_Valid_Out & channel61_Kernel17_Valid_Out & channel62_Kernel17_Valid_Out & channel63_Kernel17_Valid_Out & channel64_Kernel17_Valid_Out;

	wire channel1_Kernel18_Valid_Out, channel2_Kernel18_Valid_Out, channel3_Kernel18_Valid_Out, channel4_Kernel18_Valid_Out, channel5_Kernel18_Valid_Out, channel6_Kernel18_Valid_Out, channel7_Kernel18_Valid_Out, channel8_Kernel18_Valid_Out, channel9_Kernel18_Valid_Out, channel10_Kernel18_Valid_Out, channel11_Kernel18_Valid_Out, channel12_Kernel18_Valid_Out, channel13_Kernel18_Valid_Out, channel14_Kernel18_Valid_Out, channel15_Kernel18_Valid_Out, channel16_Kernel18_Valid_Out, channel17_Kernel18_Valid_Out, channel18_Kernel18_Valid_Out, channel19_Kernel18_Valid_Out, channel20_Kernel18_Valid_Out, channel21_Kernel18_Valid_Out, channel22_Kernel18_Valid_Out, channel23_Kernel18_Valid_Out, channel24_Kernel18_Valid_Out, channel25_Kernel18_Valid_Out, channel26_Kernel18_Valid_Out, channel27_Kernel18_Valid_Out, channel28_Kernel18_Valid_Out, channel29_Kernel18_Valid_Out, channel30_Kernel18_Valid_Out, channel31_Kernel18_Valid_Out, channel32_Kernel18_Valid_Out, channel33_Kernel18_Valid_Out, channel34_Kernel18_Valid_Out, channel35_Kernel18_Valid_Out, channel36_Kernel18_Valid_Out, channel37_Kernel18_Valid_Out, channel38_Kernel18_Valid_Out, channel39_Kernel18_Valid_Out, channel40_Kernel18_Valid_Out, channel41_Kernel18_Valid_Out, channel42_Kernel18_Valid_Out, channel43_Kernel18_Valid_Out, channel44_Kernel18_Valid_Out, channel45_Kernel18_Valid_Out, channel46_Kernel18_Valid_Out, channel47_Kernel18_Valid_Out, channel48_Kernel18_Valid_Out, channel49_Kernel18_Valid_Out, channel50_Kernel18_Valid_Out, channel51_Kernel18_Valid_Out, channel52_Kernel18_Valid_Out, channel53_Kernel18_Valid_Out, channel54_Kernel18_Valid_Out, channel55_Kernel18_Valid_Out, channel56_Kernel18_Valid_Out, channel57_Kernel18_Valid_Out, channel58_Kernel18_Valid_Out, channel59_Kernel18_Valid_Out, channel60_Kernel18_Valid_Out, channel61_Kernel18_Valid_Out, channel62_Kernel18_Valid_Out, channel63_Kernel18_Valid_Out, channel64_Kernel18_Valid_Out;

	assign add_kernel18=channel1_Kernel18_Valid_Out & channel2_Kernel18_Valid_Out & channel3_Kernel18_Valid_Out & channel4_Kernel18_Valid_Out & channel5_Kernel18_Valid_Out & channel6_Kernel18_Valid_Out & channel7_Kernel18_Valid_Out & channel8_Kernel18_Valid_Out & channel9_Kernel18_Valid_Out & channel10_Kernel18_Valid_Out & channel11_Kernel18_Valid_Out & channel12_Kernel18_Valid_Out & channel13_Kernel18_Valid_Out & channel14_Kernel18_Valid_Out & channel15_Kernel18_Valid_Out & channel16_Kernel18_Valid_Out & channel17_Kernel18_Valid_Out & channel18_Kernel18_Valid_Out & channel19_Kernel18_Valid_Out & channel20_Kernel18_Valid_Out & channel21_Kernel18_Valid_Out & channel22_Kernel18_Valid_Out & channel23_Kernel18_Valid_Out & channel24_Kernel18_Valid_Out & channel25_Kernel18_Valid_Out & channel26_Kernel18_Valid_Out & channel27_Kernel18_Valid_Out & channel28_Kernel18_Valid_Out & channel29_Kernel18_Valid_Out & channel30_Kernel18_Valid_Out & channel31_Kernel18_Valid_Out & channel32_Kernel18_Valid_Out & channel33_Kernel18_Valid_Out & channel34_Kernel18_Valid_Out & channel35_Kernel18_Valid_Out & channel36_Kernel18_Valid_Out & channel37_Kernel18_Valid_Out & channel38_Kernel18_Valid_Out & channel39_Kernel18_Valid_Out & channel40_Kernel18_Valid_Out & channel41_Kernel18_Valid_Out & channel42_Kernel18_Valid_Out & channel43_Kernel18_Valid_Out & channel44_Kernel18_Valid_Out & channel45_Kernel18_Valid_Out & channel46_Kernel18_Valid_Out & channel47_Kernel18_Valid_Out & channel48_Kernel18_Valid_Out & channel49_Kernel18_Valid_Out & channel50_Kernel18_Valid_Out & channel51_Kernel18_Valid_Out & channel52_Kernel18_Valid_Out & channel53_Kernel18_Valid_Out & channel54_Kernel18_Valid_Out & channel55_Kernel18_Valid_Out & channel56_Kernel18_Valid_Out & channel57_Kernel18_Valid_Out & channel58_Kernel18_Valid_Out & channel59_Kernel18_Valid_Out & channel60_Kernel18_Valid_Out & channel61_Kernel18_Valid_Out & channel62_Kernel18_Valid_Out & channel63_Kernel18_Valid_Out & channel64_Kernel18_Valid_Out;

	wire channel1_Kernel19_Valid_Out, channel2_Kernel19_Valid_Out, channel3_Kernel19_Valid_Out, channel4_Kernel19_Valid_Out, channel5_Kernel19_Valid_Out, channel6_Kernel19_Valid_Out, channel7_Kernel19_Valid_Out, channel8_Kernel19_Valid_Out, channel9_Kernel19_Valid_Out, channel10_Kernel19_Valid_Out, channel11_Kernel19_Valid_Out, channel12_Kernel19_Valid_Out, channel13_Kernel19_Valid_Out, channel14_Kernel19_Valid_Out, channel15_Kernel19_Valid_Out, channel16_Kernel19_Valid_Out, channel17_Kernel19_Valid_Out, channel18_Kernel19_Valid_Out, channel19_Kernel19_Valid_Out, channel20_Kernel19_Valid_Out, channel21_Kernel19_Valid_Out, channel22_Kernel19_Valid_Out, channel23_Kernel19_Valid_Out, channel24_Kernel19_Valid_Out, channel25_Kernel19_Valid_Out, channel26_Kernel19_Valid_Out, channel27_Kernel19_Valid_Out, channel28_Kernel19_Valid_Out, channel29_Kernel19_Valid_Out, channel30_Kernel19_Valid_Out, channel31_Kernel19_Valid_Out, channel32_Kernel19_Valid_Out, channel33_Kernel19_Valid_Out, channel34_Kernel19_Valid_Out, channel35_Kernel19_Valid_Out, channel36_Kernel19_Valid_Out, channel37_Kernel19_Valid_Out, channel38_Kernel19_Valid_Out, channel39_Kernel19_Valid_Out, channel40_Kernel19_Valid_Out, channel41_Kernel19_Valid_Out, channel42_Kernel19_Valid_Out, channel43_Kernel19_Valid_Out, channel44_Kernel19_Valid_Out, channel45_Kernel19_Valid_Out, channel46_Kernel19_Valid_Out, channel47_Kernel19_Valid_Out, channel48_Kernel19_Valid_Out, channel49_Kernel19_Valid_Out, channel50_Kernel19_Valid_Out, channel51_Kernel19_Valid_Out, channel52_Kernel19_Valid_Out, channel53_Kernel19_Valid_Out, channel54_Kernel19_Valid_Out, channel55_Kernel19_Valid_Out, channel56_Kernel19_Valid_Out, channel57_Kernel19_Valid_Out, channel58_Kernel19_Valid_Out, channel59_Kernel19_Valid_Out, channel60_Kernel19_Valid_Out, channel61_Kernel19_Valid_Out, channel62_Kernel19_Valid_Out, channel63_Kernel19_Valid_Out, channel64_Kernel19_Valid_Out;

	assign add_kernel19=channel1_Kernel19_Valid_Out & channel2_Kernel19_Valid_Out & channel3_Kernel19_Valid_Out & channel4_Kernel19_Valid_Out & channel5_Kernel19_Valid_Out & channel6_Kernel19_Valid_Out & channel7_Kernel19_Valid_Out & channel8_Kernel19_Valid_Out & channel9_Kernel19_Valid_Out & channel10_Kernel19_Valid_Out & channel11_Kernel19_Valid_Out & channel12_Kernel19_Valid_Out & channel13_Kernel19_Valid_Out & channel14_Kernel19_Valid_Out & channel15_Kernel19_Valid_Out & channel16_Kernel19_Valid_Out & channel17_Kernel19_Valid_Out & channel18_Kernel19_Valid_Out & channel19_Kernel19_Valid_Out & channel20_Kernel19_Valid_Out & channel21_Kernel19_Valid_Out & channel22_Kernel19_Valid_Out & channel23_Kernel19_Valid_Out & channel24_Kernel19_Valid_Out & channel25_Kernel19_Valid_Out & channel26_Kernel19_Valid_Out & channel27_Kernel19_Valid_Out & channel28_Kernel19_Valid_Out & channel29_Kernel19_Valid_Out & channel30_Kernel19_Valid_Out & channel31_Kernel19_Valid_Out & channel32_Kernel19_Valid_Out & channel33_Kernel19_Valid_Out & channel34_Kernel19_Valid_Out & channel35_Kernel19_Valid_Out & channel36_Kernel19_Valid_Out & channel37_Kernel19_Valid_Out & channel38_Kernel19_Valid_Out & channel39_Kernel19_Valid_Out & channel40_Kernel19_Valid_Out & channel41_Kernel19_Valid_Out & channel42_Kernel19_Valid_Out & channel43_Kernel19_Valid_Out & channel44_Kernel19_Valid_Out & channel45_Kernel19_Valid_Out & channel46_Kernel19_Valid_Out & channel47_Kernel19_Valid_Out & channel48_Kernel19_Valid_Out & channel49_Kernel19_Valid_Out & channel50_Kernel19_Valid_Out & channel51_Kernel19_Valid_Out & channel52_Kernel19_Valid_Out & channel53_Kernel19_Valid_Out & channel54_Kernel19_Valid_Out & channel55_Kernel19_Valid_Out & channel56_Kernel19_Valid_Out & channel57_Kernel19_Valid_Out & channel58_Kernel19_Valid_Out & channel59_Kernel19_Valid_Out & channel60_Kernel19_Valid_Out & channel61_Kernel19_Valid_Out & channel62_Kernel19_Valid_Out & channel63_Kernel19_Valid_Out & channel64_Kernel19_Valid_Out;

	wire channel1_Kernel20_Valid_Out, channel2_Kernel20_Valid_Out, channel3_Kernel20_Valid_Out, channel4_Kernel20_Valid_Out, channel5_Kernel20_Valid_Out, channel6_Kernel20_Valid_Out, channel7_Kernel20_Valid_Out, channel8_Kernel20_Valid_Out, channel9_Kernel20_Valid_Out, channel10_Kernel20_Valid_Out, channel11_Kernel20_Valid_Out, channel12_Kernel20_Valid_Out, channel13_Kernel20_Valid_Out, channel14_Kernel20_Valid_Out, channel15_Kernel20_Valid_Out, channel16_Kernel20_Valid_Out, channel17_Kernel20_Valid_Out, channel18_Kernel20_Valid_Out, channel19_Kernel20_Valid_Out, channel20_Kernel20_Valid_Out, channel21_Kernel20_Valid_Out, channel22_Kernel20_Valid_Out, channel23_Kernel20_Valid_Out, channel24_Kernel20_Valid_Out, channel25_Kernel20_Valid_Out, channel26_Kernel20_Valid_Out, channel27_Kernel20_Valid_Out, channel28_Kernel20_Valid_Out, channel29_Kernel20_Valid_Out, channel30_Kernel20_Valid_Out, channel31_Kernel20_Valid_Out, channel32_Kernel20_Valid_Out, channel33_Kernel20_Valid_Out, channel34_Kernel20_Valid_Out, channel35_Kernel20_Valid_Out, channel36_Kernel20_Valid_Out, channel37_Kernel20_Valid_Out, channel38_Kernel20_Valid_Out, channel39_Kernel20_Valid_Out, channel40_Kernel20_Valid_Out, channel41_Kernel20_Valid_Out, channel42_Kernel20_Valid_Out, channel43_Kernel20_Valid_Out, channel44_Kernel20_Valid_Out, channel45_Kernel20_Valid_Out, channel46_Kernel20_Valid_Out, channel47_Kernel20_Valid_Out, channel48_Kernel20_Valid_Out, channel49_Kernel20_Valid_Out, channel50_Kernel20_Valid_Out, channel51_Kernel20_Valid_Out, channel52_Kernel20_Valid_Out, channel53_Kernel20_Valid_Out, channel54_Kernel20_Valid_Out, channel55_Kernel20_Valid_Out, channel56_Kernel20_Valid_Out, channel57_Kernel20_Valid_Out, channel58_Kernel20_Valid_Out, channel59_Kernel20_Valid_Out, channel60_Kernel20_Valid_Out, channel61_Kernel20_Valid_Out, channel62_Kernel20_Valid_Out, channel63_Kernel20_Valid_Out, channel64_Kernel20_Valid_Out;

	assign add_kernel20=channel1_Kernel20_Valid_Out & channel2_Kernel20_Valid_Out & channel3_Kernel20_Valid_Out & channel4_Kernel20_Valid_Out & channel5_Kernel20_Valid_Out & channel6_Kernel20_Valid_Out & channel7_Kernel20_Valid_Out & channel8_Kernel20_Valid_Out & channel9_Kernel20_Valid_Out & channel10_Kernel20_Valid_Out & channel11_Kernel20_Valid_Out & channel12_Kernel20_Valid_Out & channel13_Kernel20_Valid_Out & channel14_Kernel20_Valid_Out & channel15_Kernel20_Valid_Out & channel16_Kernel20_Valid_Out & channel17_Kernel20_Valid_Out & channel18_Kernel20_Valid_Out & channel19_Kernel20_Valid_Out & channel20_Kernel20_Valid_Out & channel21_Kernel20_Valid_Out & channel22_Kernel20_Valid_Out & channel23_Kernel20_Valid_Out & channel24_Kernel20_Valid_Out & channel25_Kernel20_Valid_Out & channel26_Kernel20_Valid_Out & channel27_Kernel20_Valid_Out & channel28_Kernel20_Valid_Out & channel29_Kernel20_Valid_Out & channel30_Kernel20_Valid_Out & channel31_Kernel20_Valid_Out & channel32_Kernel20_Valid_Out & channel33_Kernel20_Valid_Out & channel34_Kernel20_Valid_Out & channel35_Kernel20_Valid_Out & channel36_Kernel20_Valid_Out & channel37_Kernel20_Valid_Out & channel38_Kernel20_Valid_Out & channel39_Kernel20_Valid_Out & channel40_Kernel20_Valid_Out & channel41_Kernel20_Valid_Out & channel42_Kernel20_Valid_Out & channel43_Kernel20_Valid_Out & channel44_Kernel20_Valid_Out & channel45_Kernel20_Valid_Out & channel46_Kernel20_Valid_Out & channel47_Kernel20_Valid_Out & channel48_Kernel20_Valid_Out & channel49_Kernel20_Valid_Out & channel50_Kernel20_Valid_Out & channel51_Kernel20_Valid_Out & channel52_Kernel20_Valid_Out & channel53_Kernel20_Valid_Out & channel54_Kernel20_Valid_Out & channel55_Kernel20_Valid_Out & channel56_Kernel20_Valid_Out & channel57_Kernel20_Valid_Out & channel58_Kernel20_Valid_Out & channel59_Kernel20_Valid_Out & channel60_Kernel20_Valid_Out & channel61_Kernel20_Valid_Out & channel62_Kernel20_Valid_Out & channel63_Kernel20_Valid_Out & channel64_Kernel20_Valid_Out;

	wire channel1_Kernel21_Valid_Out, channel2_Kernel21_Valid_Out, channel3_Kernel21_Valid_Out, channel4_Kernel21_Valid_Out, channel5_Kernel21_Valid_Out, channel6_Kernel21_Valid_Out, channel7_Kernel21_Valid_Out, channel8_Kernel21_Valid_Out, channel9_Kernel21_Valid_Out, channel10_Kernel21_Valid_Out, channel11_Kernel21_Valid_Out, channel12_Kernel21_Valid_Out, channel13_Kernel21_Valid_Out, channel14_Kernel21_Valid_Out, channel15_Kernel21_Valid_Out, channel16_Kernel21_Valid_Out, channel17_Kernel21_Valid_Out, channel18_Kernel21_Valid_Out, channel19_Kernel21_Valid_Out, channel20_Kernel21_Valid_Out, channel21_Kernel21_Valid_Out, channel22_Kernel21_Valid_Out, channel23_Kernel21_Valid_Out, channel24_Kernel21_Valid_Out, channel25_Kernel21_Valid_Out, channel26_Kernel21_Valid_Out, channel27_Kernel21_Valid_Out, channel28_Kernel21_Valid_Out, channel29_Kernel21_Valid_Out, channel30_Kernel21_Valid_Out, channel31_Kernel21_Valid_Out, channel32_Kernel21_Valid_Out, channel33_Kernel21_Valid_Out, channel34_Kernel21_Valid_Out, channel35_Kernel21_Valid_Out, channel36_Kernel21_Valid_Out, channel37_Kernel21_Valid_Out, channel38_Kernel21_Valid_Out, channel39_Kernel21_Valid_Out, channel40_Kernel21_Valid_Out, channel41_Kernel21_Valid_Out, channel42_Kernel21_Valid_Out, channel43_Kernel21_Valid_Out, channel44_Kernel21_Valid_Out, channel45_Kernel21_Valid_Out, channel46_Kernel21_Valid_Out, channel47_Kernel21_Valid_Out, channel48_Kernel21_Valid_Out, channel49_Kernel21_Valid_Out, channel50_Kernel21_Valid_Out, channel51_Kernel21_Valid_Out, channel52_Kernel21_Valid_Out, channel53_Kernel21_Valid_Out, channel54_Kernel21_Valid_Out, channel55_Kernel21_Valid_Out, channel56_Kernel21_Valid_Out, channel57_Kernel21_Valid_Out, channel58_Kernel21_Valid_Out, channel59_Kernel21_Valid_Out, channel60_Kernel21_Valid_Out, channel61_Kernel21_Valid_Out, channel62_Kernel21_Valid_Out, channel63_Kernel21_Valid_Out, channel64_Kernel21_Valid_Out;

	assign add_kernel21=channel1_Kernel21_Valid_Out & channel2_Kernel21_Valid_Out & channel3_Kernel21_Valid_Out & channel4_Kernel21_Valid_Out & channel5_Kernel21_Valid_Out & channel6_Kernel21_Valid_Out & channel7_Kernel21_Valid_Out & channel8_Kernel21_Valid_Out & channel9_Kernel21_Valid_Out & channel10_Kernel21_Valid_Out & channel11_Kernel21_Valid_Out & channel12_Kernel21_Valid_Out & channel13_Kernel21_Valid_Out & channel14_Kernel21_Valid_Out & channel15_Kernel21_Valid_Out & channel16_Kernel21_Valid_Out & channel17_Kernel21_Valid_Out & channel18_Kernel21_Valid_Out & channel19_Kernel21_Valid_Out & channel20_Kernel21_Valid_Out & channel21_Kernel21_Valid_Out & channel22_Kernel21_Valid_Out & channel23_Kernel21_Valid_Out & channel24_Kernel21_Valid_Out & channel25_Kernel21_Valid_Out & channel26_Kernel21_Valid_Out & channel27_Kernel21_Valid_Out & channel28_Kernel21_Valid_Out & channel29_Kernel21_Valid_Out & channel30_Kernel21_Valid_Out & channel31_Kernel21_Valid_Out & channel32_Kernel21_Valid_Out & channel33_Kernel21_Valid_Out & channel34_Kernel21_Valid_Out & channel35_Kernel21_Valid_Out & channel36_Kernel21_Valid_Out & channel37_Kernel21_Valid_Out & channel38_Kernel21_Valid_Out & channel39_Kernel21_Valid_Out & channel40_Kernel21_Valid_Out & channel41_Kernel21_Valid_Out & channel42_Kernel21_Valid_Out & channel43_Kernel21_Valid_Out & channel44_Kernel21_Valid_Out & channel45_Kernel21_Valid_Out & channel46_Kernel21_Valid_Out & channel47_Kernel21_Valid_Out & channel48_Kernel21_Valid_Out & channel49_Kernel21_Valid_Out & channel50_Kernel21_Valid_Out & channel51_Kernel21_Valid_Out & channel52_Kernel21_Valid_Out & channel53_Kernel21_Valid_Out & channel54_Kernel21_Valid_Out & channel55_Kernel21_Valid_Out & channel56_Kernel21_Valid_Out & channel57_Kernel21_Valid_Out & channel58_Kernel21_Valid_Out & channel59_Kernel21_Valid_Out & channel60_Kernel21_Valid_Out & channel61_Kernel21_Valid_Out & channel62_Kernel21_Valid_Out & channel63_Kernel21_Valid_Out & channel64_Kernel21_Valid_Out;

	wire channel1_Kernel22_Valid_Out, channel2_Kernel22_Valid_Out, channel3_Kernel22_Valid_Out, channel4_Kernel22_Valid_Out, channel5_Kernel22_Valid_Out, channel6_Kernel22_Valid_Out, channel7_Kernel22_Valid_Out, channel8_Kernel22_Valid_Out, channel9_Kernel22_Valid_Out, channel10_Kernel22_Valid_Out, channel11_Kernel22_Valid_Out, channel12_Kernel22_Valid_Out, channel13_Kernel22_Valid_Out, channel14_Kernel22_Valid_Out, channel15_Kernel22_Valid_Out, channel16_Kernel22_Valid_Out, channel17_Kernel22_Valid_Out, channel18_Kernel22_Valid_Out, channel19_Kernel22_Valid_Out, channel20_Kernel22_Valid_Out, channel21_Kernel22_Valid_Out, channel22_Kernel22_Valid_Out, channel23_Kernel22_Valid_Out, channel24_Kernel22_Valid_Out, channel25_Kernel22_Valid_Out, channel26_Kernel22_Valid_Out, channel27_Kernel22_Valid_Out, channel28_Kernel22_Valid_Out, channel29_Kernel22_Valid_Out, channel30_Kernel22_Valid_Out, channel31_Kernel22_Valid_Out, channel32_Kernel22_Valid_Out, channel33_Kernel22_Valid_Out, channel34_Kernel22_Valid_Out, channel35_Kernel22_Valid_Out, channel36_Kernel22_Valid_Out, channel37_Kernel22_Valid_Out, channel38_Kernel22_Valid_Out, channel39_Kernel22_Valid_Out, channel40_Kernel22_Valid_Out, channel41_Kernel22_Valid_Out, channel42_Kernel22_Valid_Out, channel43_Kernel22_Valid_Out, channel44_Kernel22_Valid_Out, channel45_Kernel22_Valid_Out, channel46_Kernel22_Valid_Out, channel47_Kernel22_Valid_Out, channel48_Kernel22_Valid_Out, channel49_Kernel22_Valid_Out, channel50_Kernel22_Valid_Out, channel51_Kernel22_Valid_Out, channel52_Kernel22_Valid_Out, channel53_Kernel22_Valid_Out, channel54_Kernel22_Valid_Out, channel55_Kernel22_Valid_Out, channel56_Kernel22_Valid_Out, channel57_Kernel22_Valid_Out, channel58_Kernel22_Valid_Out, channel59_Kernel22_Valid_Out, channel60_Kernel22_Valid_Out, channel61_Kernel22_Valid_Out, channel62_Kernel22_Valid_Out, channel63_Kernel22_Valid_Out, channel64_Kernel22_Valid_Out;

	assign add_kernel22=channel1_Kernel22_Valid_Out & channel2_Kernel22_Valid_Out & channel3_Kernel22_Valid_Out & channel4_Kernel22_Valid_Out & channel5_Kernel22_Valid_Out & channel6_Kernel22_Valid_Out & channel7_Kernel22_Valid_Out & channel8_Kernel22_Valid_Out & channel9_Kernel22_Valid_Out & channel10_Kernel22_Valid_Out & channel11_Kernel22_Valid_Out & channel12_Kernel22_Valid_Out & channel13_Kernel22_Valid_Out & channel14_Kernel22_Valid_Out & channel15_Kernel22_Valid_Out & channel16_Kernel22_Valid_Out & channel17_Kernel22_Valid_Out & channel18_Kernel22_Valid_Out & channel19_Kernel22_Valid_Out & channel20_Kernel22_Valid_Out & channel21_Kernel22_Valid_Out & channel22_Kernel22_Valid_Out & channel23_Kernel22_Valid_Out & channel24_Kernel22_Valid_Out & channel25_Kernel22_Valid_Out & channel26_Kernel22_Valid_Out & channel27_Kernel22_Valid_Out & channel28_Kernel22_Valid_Out & channel29_Kernel22_Valid_Out & channel30_Kernel22_Valid_Out & channel31_Kernel22_Valid_Out & channel32_Kernel22_Valid_Out & channel33_Kernel22_Valid_Out & channel34_Kernel22_Valid_Out & channel35_Kernel22_Valid_Out & channel36_Kernel22_Valid_Out & channel37_Kernel22_Valid_Out & channel38_Kernel22_Valid_Out & channel39_Kernel22_Valid_Out & channel40_Kernel22_Valid_Out & channel41_Kernel22_Valid_Out & channel42_Kernel22_Valid_Out & channel43_Kernel22_Valid_Out & channel44_Kernel22_Valid_Out & channel45_Kernel22_Valid_Out & channel46_Kernel22_Valid_Out & channel47_Kernel22_Valid_Out & channel48_Kernel22_Valid_Out & channel49_Kernel22_Valid_Out & channel50_Kernel22_Valid_Out & channel51_Kernel22_Valid_Out & channel52_Kernel22_Valid_Out & channel53_Kernel22_Valid_Out & channel54_Kernel22_Valid_Out & channel55_Kernel22_Valid_Out & channel56_Kernel22_Valid_Out & channel57_Kernel22_Valid_Out & channel58_Kernel22_Valid_Out & channel59_Kernel22_Valid_Out & channel60_Kernel22_Valid_Out & channel61_Kernel22_Valid_Out & channel62_Kernel22_Valid_Out & channel63_Kernel22_Valid_Out & channel64_Kernel22_Valid_Out;

	wire channel1_Kernel23_Valid_Out, channel2_Kernel23_Valid_Out, channel3_Kernel23_Valid_Out, channel4_Kernel23_Valid_Out, channel5_Kernel23_Valid_Out, channel6_Kernel23_Valid_Out, channel7_Kernel23_Valid_Out, channel8_Kernel23_Valid_Out, channel9_Kernel23_Valid_Out, channel10_Kernel23_Valid_Out, channel11_Kernel23_Valid_Out, channel12_Kernel23_Valid_Out, channel13_Kernel23_Valid_Out, channel14_Kernel23_Valid_Out, channel15_Kernel23_Valid_Out, channel16_Kernel23_Valid_Out, channel17_Kernel23_Valid_Out, channel18_Kernel23_Valid_Out, channel19_Kernel23_Valid_Out, channel20_Kernel23_Valid_Out, channel21_Kernel23_Valid_Out, channel22_Kernel23_Valid_Out, channel23_Kernel23_Valid_Out, channel24_Kernel23_Valid_Out, channel25_Kernel23_Valid_Out, channel26_Kernel23_Valid_Out, channel27_Kernel23_Valid_Out, channel28_Kernel23_Valid_Out, channel29_Kernel23_Valid_Out, channel30_Kernel23_Valid_Out, channel31_Kernel23_Valid_Out, channel32_Kernel23_Valid_Out, channel33_Kernel23_Valid_Out, channel34_Kernel23_Valid_Out, channel35_Kernel23_Valid_Out, channel36_Kernel23_Valid_Out, channel37_Kernel23_Valid_Out, channel38_Kernel23_Valid_Out, channel39_Kernel23_Valid_Out, channel40_Kernel23_Valid_Out, channel41_Kernel23_Valid_Out, channel42_Kernel23_Valid_Out, channel43_Kernel23_Valid_Out, channel44_Kernel23_Valid_Out, channel45_Kernel23_Valid_Out, channel46_Kernel23_Valid_Out, channel47_Kernel23_Valid_Out, channel48_Kernel23_Valid_Out, channel49_Kernel23_Valid_Out, channel50_Kernel23_Valid_Out, channel51_Kernel23_Valid_Out, channel52_Kernel23_Valid_Out, channel53_Kernel23_Valid_Out, channel54_Kernel23_Valid_Out, channel55_Kernel23_Valid_Out, channel56_Kernel23_Valid_Out, channel57_Kernel23_Valid_Out, channel58_Kernel23_Valid_Out, channel59_Kernel23_Valid_Out, channel60_Kernel23_Valid_Out, channel61_Kernel23_Valid_Out, channel62_Kernel23_Valid_Out, channel63_Kernel23_Valid_Out, channel64_Kernel23_Valid_Out;

	assign add_kernel23=channel1_Kernel23_Valid_Out & channel2_Kernel23_Valid_Out & channel3_Kernel23_Valid_Out & channel4_Kernel23_Valid_Out & channel5_Kernel23_Valid_Out & channel6_Kernel23_Valid_Out & channel7_Kernel23_Valid_Out & channel8_Kernel23_Valid_Out & channel9_Kernel23_Valid_Out & channel10_Kernel23_Valid_Out & channel11_Kernel23_Valid_Out & channel12_Kernel23_Valid_Out & channel13_Kernel23_Valid_Out & channel14_Kernel23_Valid_Out & channel15_Kernel23_Valid_Out & channel16_Kernel23_Valid_Out & channel17_Kernel23_Valid_Out & channel18_Kernel23_Valid_Out & channel19_Kernel23_Valid_Out & channel20_Kernel23_Valid_Out & channel21_Kernel23_Valid_Out & channel22_Kernel23_Valid_Out & channel23_Kernel23_Valid_Out & channel24_Kernel23_Valid_Out & channel25_Kernel23_Valid_Out & channel26_Kernel23_Valid_Out & channel27_Kernel23_Valid_Out & channel28_Kernel23_Valid_Out & channel29_Kernel23_Valid_Out & channel30_Kernel23_Valid_Out & channel31_Kernel23_Valid_Out & channel32_Kernel23_Valid_Out & channel33_Kernel23_Valid_Out & channel34_Kernel23_Valid_Out & channel35_Kernel23_Valid_Out & channel36_Kernel23_Valid_Out & channel37_Kernel23_Valid_Out & channel38_Kernel23_Valid_Out & channel39_Kernel23_Valid_Out & channel40_Kernel23_Valid_Out & channel41_Kernel23_Valid_Out & channel42_Kernel23_Valid_Out & channel43_Kernel23_Valid_Out & channel44_Kernel23_Valid_Out & channel45_Kernel23_Valid_Out & channel46_Kernel23_Valid_Out & channel47_Kernel23_Valid_Out & channel48_Kernel23_Valid_Out & channel49_Kernel23_Valid_Out & channel50_Kernel23_Valid_Out & channel51_Kernel23_Valid_Out & channel52_Kernel23_Valid_Out & channel53_Kernel23_Valid_Out & channel54_Kernel23_Valid_Out & channel55_Kernel23_Valid_Out & channel56_Kernel23_Valid_Out & channel57_Kernel23_Valid_Out & channel58_Kernel23_Valid_Out & channel59_Kernel23_Valid_Out & channel60_Kernel23_Valid_Out & channel61_Kernel23_Valid_Out & channel62_Kernel23_Valid_Out & channel63_Kernel23_Valid_Out & channel64_Kernel23_Valid_Out;

	wire channel1_Kernel24_Valid_Out, channel2_Kernel24_Valid_Out, channel3_Kernel24_Valid_Out, channel4_Kernel24_Valid_Out, channel5_Kernel24_Valid_Out, channel6_Kernel24_Valid_Out, channel7_Kernel24_Valid_Out, channel8_Kernel24_Valid_Out, channel9_Kernel24_Valid_Out, channel10_Kernel24_Valid_Out, channel11_Kernel24_Valid_Out, channel12_Kernel24_Valid_Out, channel13_Kernel24_Valid_Out, channel14_Kernel24_Valid_Out, channel15_Kernel24_Valid_Out, channel16_Kernel24_Valid_Out, channel17_Kernel24_Valid_Out, channel18_Kernel24_Valid_Out, channel19_Kernel24_Valid_Out, channel20_Kernel24_Valid_Out, channel21_Kernel24_Valid_Out, channel22_Kernel24_Valid_Out, channel23_Kernel24_Valid_Out, channel24_Kernel24_Valid_Out, channel25_Kernel24_Valid_Out, channel26_Kernel24_Valid_Out, channel27_Kernel24_Valid_Out, channel28_Kernel24_Valid_Out, channel29_Kernel24_Valid_Out, channel30_Kernel24_Valid_Out, channel31_Kernel24_Valid_Out, channel32_Kernel24_Valid_Out, channel33_Kernel24_Valid_Out, channel34_Kernel24_Valid_Out, channel35_Kernel24_Valid_Out, channel36_Kernel24_Valid_Out, channel37_Kernel24_Valid_Out, channel38_Kernel24_Valid_Out, channel39_Kernel24_Valid_Out, channel40_Kernel24_Valid_Out, channel41_Kernel24_Valid_Out, channel42_Kernel24_Valid_Out, channel43_Kernel24_Valid_Out, channel44_Kernel24_Valid_Out, channel45_Kernel24_Valid_Out, channel46_Kernel24_Valid_Out, channel47_Kernel24_Valid_Out, channel48_Kernel24_Valid_Out, channel49_Kernel24_Valid_Out, channel50_Kernel24_Valid_Out, channel51_Kernel24_Valid_Out, channel52_Kernel24_Valid_Out, channel53_Kernel24_Valid_Out, channel54_Kernel24_Valid_Out, channel55_Kernel24_Valid_Out, channel56_Kernel24_Valid_Out, channel57_Kernel24_Valid_Out, channel58_Kernel24_Valid_Out, channel59_Kernel24_Valid_Out, channel60_Kernel24_Valid_Out, channel61_Kernel24_Valid_Out, channel62_Kernel24_Valid_Out, channel63_Kernel24_Valid_Out, channel64_Kernel24_Valid_Out;

	assign add_kernel24=channel1_Kernel24_Valid_Out & channel2_Kernel24_Valid_Out & channel3_Kernel24_Valid_Out & channel4_Kernel24_Valid_Out & channel5_Kernel24_Valid_Out & channel6_Kernel24_Valid_Out & channel7_Kernel24_Valid_Out & channel8_Kernel24_Valid_Out & channel9_Kernel24_Valid_Out & channel10_Kernel24_Valid_Out & channel11_Kernel24_Valid_Out & channel12_Kernel24_Valid_Out & channel13_Kernel24_Valid_Out & channel14_Kernel24_Valid_Out & channel15_Kernel24_Valid_Out & channel16_Kernel24_Valid_Out & channel17_Kernel24_Valid_Out & channel18_Kernel24_Valid_Out & channel19_Kernel24_Valid_Out & channel20_Kernel24_Valid_Out & channel21_Kernel24_Valid_Out & channel22_Kernel24_Valid_Out & channel23_Kernel24_Valid_Out & channel24_Kernel24_Valid_Out & channel25_Kernel24_Valid_Out & channel26_Kernel24_Valid_Out & channel27_Kernel24_Valid_Out & channel28_Kernel24_Valid_Out & channel29_Kernel24_Valid_Out & channel30_Kernel24_Valid_Out & channel31_Kernel24_Valid_Out & channel32_Kernel24_Valid_Out & channel33_Kernel24_Valid_Out & channel34_Kernel24_Valid_Out & channel35_Kernel24_Valid_Out & channel36_Kernel24_Valid_Out & channel37_Kernel24_Valid_Out & channel38_Kernel24_Valid_Out & channel39_Kernel24_Valid_Out & channel40_Kernel24_Valid_Out & channel41_Kernel24_Valid_Out & channel42_Kernel24_Valid_Out & channel43_Kernel24_Valid_Out & channel44_Kernel24_Valid_Out & channel45_Kernel24_Valid_Out & channel46_Kernel24_Valid_Out & channel47_Kernel24_Valid_Out & channel48_Kernel24_Valid_Out & channel49_Kernel24_Valid_Out & channel50_Kernel24_Valid_Out & channel51_Kernel24_Valid_Out & channel52_Kernel24_Valid_Out & channel53_Kernel24_Valid_Out & channel54_Kernel24_Valid_Out & channel55_Kernel24_Valid_Out & channel56_Kernel24_Valid_Out & channel57_Kernel24_Valid_Out & channel58_Kernel24_Valid_Out & channel59_Kernel24_Valid_Out & channel60_Kernel24_Valid_Out & channel61_Kernel24_Valid_Out & channel62_Kernel24_Valid_Out & channel63_Kernel24_Valid_Out & channel64_Kernel24_Valid_Out;

	wire channel1_Kernel25_Valid_Out, channel2_Kernel25_Valid_Out, channel3_Kernel25_Valid_Out, channel4_Kernel25_Valid_Out, channel5_Kernel25_Valid_Out, channel6_Kernel25_Valid_Out, channel7_Kernel25_Valid_Out, channel8_Kernel25_Valid_Out, channel9_Kernel25_Valid_Out, channel10_Kernel25_Valid_Out, channel11_Kernel25_Valid_Out, channel12_Kernel25_Valid_Out, channel13_Kernel25_Valid_Out, channel14_Kernel25_Valid_Out, channel15_Kernel25_Valid_Out, channel16_Kernel25_Valid_Out, channel17_Kernel25_Valid_Out, channel18_Kernel25_Valid_Out, channel19_Kernel25_Valid_Out, channel20_Kernel25_Valid_Out, channel21_Kernel25_Valid_Out, channel22_Kernel25_Valid_Out, channel23_Kernel25_Valid_Out, channel24_Kernel25_Valid_Out, channel25_Kernel25_Valid_Out, channel26_Kernel25_Valid_Out, channel27_Kernel25_Valid_Out, channel28_Kernel25_Valid_Out, channel29_Kernel25_Valid_Out, channel30_Kernel25_Valid_Out, channel31_Kernel25_Valid_Out, channel32_Kernel25_Valid_Out, channel33_Kernel25_Valid_Out, channel34_Kernel25_Valid_Out, channel35_Kernel25_Valid_Out, channel36_Kernel25_Valid_Out, channel37_Kernel25_Valid_Out, channel38_Kernel25_Valid_Out, channel39_Kernel25_Valid_Out, channel40_Kernel25_Valid_Out, channel41_Kernel25_Valid_Out, channel42_Kernel25_Valid_Out, channel43_Kernel25_Valid_Out, channel44_Kernel25_Valid_Out, channel45_Kernel25_Valid_Out, channel46_Kernel25_Valid_Out, channel47_Kernel25_Valid_Out, channel48_Kernel25_Valid_Out, channel49_Kernel25_Valid_Out, channel50_Kernel25_Valid_Out, channel51_Kernel25_Valid_Out, channel52_Kernel25_Valid_Out, channel53_Kernel25_Valid_Out, channel54_Kernel25_Valid_Out, channel55_Kernel25_Valid_Out, channel56_Kernel25_Valid_Out, channel57_Kernel25_Valid_Out, channel58_Kernel25_Valid_Out, channel59_Kernel25_Valid_Out, channel60_Kernel25_Valid_Out, channel61_Kernel25_Valid_Out, channel62_Kernel25_Valid_Out, channel63_Kernel25_Valid_Out, channel64_Kernel25_Valid_Out;

	assign add_kernel25=channel1_Kernel25_Valid_Out & channel2_Kernel25_Valid_Out & channel3_Kernel25_Valid_Out & channel4_Kernel25_Valid_Out & channel5_Kernel25_Valid_Out & channel6_Kernel25_Valid_Out & channel7_Kernel25_Valid_Out & channel8_Kernel25_Valid_Out & channel9_Kernel25_Valid_Out & channel10_Kernel25_Valid_Out & channel11_Kernel25_Valid_Out & channel12_Kernel25_Valid_Out & channel13_Kernel25_Valid_Out & channel14_Kernel25_Valid_Out & channel15_Kernel25_Valid_Out & channel16_Kernel25_Valid_Out & channel17_Kernel25_Valid_Out & channel18_Kernel25_Valid_Out & channel19_Kernel25_Valid_Out & channel20_Kernel25_Valid_Out & channel21_Kernel25_Valid_Out & channel22_Kernel25_Valid_Out & channel23_Kernel25_Valid_Out & channel24_Kernel25_Valid_Out & channel25_Kernel25_Valid_Out & channel26_Kernel25_Valid_Out & channel27_Kernel25_Valid_Out & channel28_Kernel25_Valid_Out & channel29_Kernel25_Valid_Out & channel30_Kernel25_Valid_Out & channel31_Kernel25_Valid_Out & channel32_Kernel25_Valid_Out & channel33_Kernel25_Valid_Out & channel34_Kernel25_Valid_Out & channel35_Kernel25_Valid_Out & channel36_Kernel25_Valid_Out & channel37_Kernel25_Valid_Out & channel38_Kernel25_Valid_Out & channel39_Kernel25_Valid_Out & channel40_Kernel25_Valid_Out & channel41_Kernel25_Valid_Out & channel42_Kernel25_Valid_Out & channel43_Kernel25_Valid_Out & channel44_Kernel25_Valid_Out & channel45_Kernel25_Valid_Out & channel46_Kernel25_Valid_Out & channel47_Kernel25_Valid_Out & channel48_Kernel25_Valid_Out & channel49_Kernel25_Valid_Out & channel50_Kernel25_Valid_Out & channel51_Kernel25_Valid_Out & channel52_Kernel25_Valid_Out & channel53_Kernel25_Valid_Out & channel54_Kernel25_Valid_Out & channel55_Kernel25_Valid_Out & channel56_Kernel25_Valid_Out & channel57_Kernel25_Valid_Out & channel58_Kernel25_Valid_Out & channel59_Kernel25_Valid_Out & channel60_Kernel25_Valid_Out & channel61_Kernel25_Valid_Out & channel62_Kernel25_Valid_Out & channel63_Kernel25_Valid_Out & channel64_Kernel25_Valid_Out;

	wire channel1_Kernel26_Valid_Out, channel2_Kernel26_Valid_Out, channel3_Kernel26_Valid_Out, channel4_Kernel26_Valid_Out, channel5_Kernel26_Valid_Out, channel6_Kernel26_Valid_Out, channel7_Kernel26_Valid_Out, channel8_Kernel26_Valid_Out, channel9_Kernel26_Valid_Out, channel10_Kernel26_Valid_Out, channel11_Kernel26_Valid_Out, channel12_Kernel26_Valid_Out, channel13_Kernel26_Valid_Out, channel14_Kernel26_Valid_Out, channel15_Kernel26_Valid_Out, channel16_Kernel26_Valid_Out, channel17_Kernel26_Valid_Out, channel18_Kernel26_Valid_Out, channel19_Kernel26_Valid_Out, channel20_Kernel26_Valid_Out, channel21_Kernel26_Valid_Out, channel22_Kernel26_Valid_Out, channel23_Kernel26_Valid_Out, channel24_Kernel26_Valid_Out, channel25_Kernel26_Valid_Out, channel26_Kernel26_Valid_Out, channel27_Kernel26_Valid_Out, channel28_Kernel26_Valid_Out, channel29_Kernel26_Valid_Out, channel30_Kernel26_Valid_Out, channel31_Kernel26_Valid_Out, channel32_Kernel26_Valid_Out, channel33_Kernel26_Valid_Out, channel34_Kernel26_Valid_Out, channel35_Kernel26_Valid_Out, channel36_Kernel26_Valid_Out, channel37_Kernel26_Valid_Out, channel38_Kernel26_Valid_Out, channel39_Kernel26_Valid_Out, channel40_Kernel26_Valid_Out, channel41_Kernel26_Valid_Out, channel42_Kernel26_Valid_Out, channel43_Kernel26_Valid_Out, channel44_Kernel26_Valid_Out, channel45_Kernel26_Valid_Out, channel46_Kernel26_Valid_Out, channel47_Kernel26_Valid_Out, channel48_Kernel26_Valid_Out, channel49_Kernel26_Valid_Out, channel50_Kernel26_Valid_Out, channel51_Kernel26_Valid_Out, channel52_Kernel26_Valid_Out, channel53_Kernel26_Valid_Out, channel54_Kernel26_Valid_Out, channel55_Kernel26_Valid_Out, channel56_Kernel26_Valid_Out, channel57_Kernel26_Valid_Out, channel58_Kernel26_Valid_Out, channel59_Kernel26_Valid_Out, channel60_Kernel26_Valid_Out, channel61_Kernel26_Valid_Out, channel62_Kernel26_Valid_Out, channel63_Kernel26_Valid_Out, channel64_Kernel26_Valid_Out;

	assign add_kernel26=channel1_Kernel26_Valid_Out & channel2_Kernel26_Valid_Out & channel3_Kernel26_Valid_Out & channel4_Kernel26_Valid_Out & channel5_Kernel26_Valid_Out & channel6_Kernel26_Valid_Out & channel7_Kernel26_Valid_Out & channel8_Kernel26_Valid_Out & channel9_Kernel26_Valid_Out & channel10_Kernel26_Valid_Out & channel11_Kernel26_Valid_Out & channel12_Kernel26_Valid_Out & channel13_Kernel26_Valid_Out & channel14_Kernel26_Valid_Out & channel15_Kernel26_Valid_Out & channel16_Kernel26_Valid_Out & channel17_Kernel26_Valid_Out & channel18_Kernel26_Valid_Out & channel19_Kernel26_Valid_Out & channel20_Kernel26_Valid_Out & channel21_Kernel26_Valid_Out & channel22_Kernel26_Valid_Out & channel23_Kernel26_Valid_Out & channel24_Kernel26_Valid_Out & channel25_Kernel26_Valid_Out & channel26_Kernel26_Valid_Out & channel27_Kernel26_Valid_Out & channel28_Kernel26_Valid_Out & channel29_Kernel26_Valid_Out & channel30_Kernel26_Valid_Out & channel31_Kernel26_Valid_Out & channel32_Kernel26_Valid_Out & channel33_Kernel26_Valid_Out & channel34_Kernel26_Valid_Out & channel35_Kernel26_Valid_Out & channel36_Kernel26_Valid_Out & channel37_Kernel26_Valid_Out & channel38_Kernel26_Valid_Out & channel39_Kernel26_Valid_Out & channel40_Kernel26_Valid_Out & channel41_Kernel26_Valid_Out & channel42_Kernel26_Valid_Out & channel43_Kernel26_Valid_Out & channel44_Kernel26_Valid_Out & channel45_Kernel26_Valid_Out & channel46_Kernel26_Valid_Out & channel47_Kernel26_Valid_Out & channel48_Kernel26_Valid_Out & channel49_Kernel26_Valid_Out & channel50_Kernel26_Valid_Out & channel51_Kernel26_Valid_Out & channel52_Kernel26_Valid_Out & channel53_Kernel26_Valid_Out & channel54_Kernel26_Valid_Out & channel55_Kernel26_Valid_Out & channel56_Kernel26_Valid_Out & channel57_Kernel26_Valid_Out & channel58_Kernel26_Valid_Out & channel59_Kernel26_Valid_Out & channel60_Kernel26_Valid_Out & channel61_Kernel26_Valid_Out & channel62_Kernel26_Valid_Out & channel63_Kernel26_Valid_Out & channel64_Kernel26_Valid_Out;

	wire channel1_Kernel27_Valid_Out, channel2_Kernel27_Valid_Out, channel3_Kernel27_Valid_Out, channel4_Kernel27_Valid_Out, channel5_Kernel27_Valid_Out, channel6_Kernel27_Valid_Out, channel7_Kernel27_Valid_Out, channel8_Kernel27_Valid_Out, channel9_Kernel27_Valid_Out, channel10_Kernel27_Valid_Out, channel11_Kernel27_Valid_Out, channel12_Kernel27_Valid_Out, channel13_Kernel27_Valid_Out, channel14_Kernel27_Valid_Out, channel15_Kernel27_Valid_Out, channel16_Kernel27_Valid_Out, channel17_Kernel27_Valid_Out, channel18_Kernel27_Valid_Out, channel19_Kernel27_Valid_Out, channel20_Kernel27_Valid_Out, channel21_Kernel27_Valid_Out, channel22_Kernel27_Valid_Out, channel23_Kernel27_Valid_Out, channel24_Kernel27_Valid_Out, channel25_Kernel27_Valid_Out, channel26_Kernel27_Valid_Out, channel27_Kernel27_Valid_Out, channel28_Kernel27_Valid_Out, channel29_Kernel27_Valid_Out, channel30_Kernel27_Valid_Out, channel31_Kernel27_Valid_Out, channel32_Kernel27_Valid_Out, channel33_Kernel27_Valid_Out, channel34_Kernel27_Valid_Out, channel35_Kernel27_Valid_Out, channel36_Kernel27_Valid_Out, channel37_Kernel27_Valid_Out, channel38_Kernel27_Valid_Out, channel39_Kernel27_Valid_Out, channel40_Kernel27_Valid_Out, channel41_Kernel27_Valid_Out, channel42_Kernel27_Valid_Out, channel43_Kernel27_Valid_Out, channel44_Kernel27_Valid_Out, channel45_Kernel27_Valid_Out, channel46_Kernel27_Valid_Out, channel47_Kernel27_Valid_Out, channel48_Kernel27_Valid_Out, channel49_Kernel27_Valid_Out, channel50_Kernel27_Valid_Out, channel51_Kernel27_Valid_Out, channel52_Kernel27_Valid_Out, channel53_Kernel27_Valid_Out, channel54_Kernel27_Valid_Out, channel55_Kernel27_Valid_Out, channel56_Kernel27_Valid_Out, channel57_Kernel27_Valid_Out, channel58_Kernel27_Valid_Out, channel59_Kernel27_Valid_Out, channel60_Kernel27_Valid_Out, channel61_Kernel27_Valid_Out, channel62_Kernel27_Valid_Out, channel63_Kernel27_Valid_Out, channel64_Kernel27_Valid_Out;

	assign add_kernel27=channel1_Kernel27_Valid_Out & channel2_Kernel27_Valid_Out & channel3_Kernel27_Valid_Out & channel4_Kernel27_Valid_Out & channel5_Kernel27_Valid_Out & channel6_Kernel27_Valid_Out & channel7_Kernel27_Valid_Out & channel8_Kernel27_Valid_Out & channel9_Kernel27_Valid_Out & channel10_Kernel27_Valid_Out & channel11_Kernel27_Valid_Out & channel12_Kernel27_Valid_Out & channel13_Kernel27_Valid_Out & channel14_Kernel27_Valid_Out & channel15_Kernel27_Valid_Out & channel16_Kernel27_Valid_Out & channel17_Kernel27_Valid_Out & channel18_Kernel27_Valid_Out & channel19_Kernel27_Valid_Out & channel20_Kernel27_Valid_Out & channel21_Kernel27_Valid_Out & channel22_Kernel27_Valid_Out & channel23_Kernel27_Valid_Out & channel24_Kernel27_Valid_Out & channel25_Kernel27_Valid_Out & channel26_Kernel27_Valid_Out & channel27_Kernel27_Valid_Out & channel28_Kernel27_Valid_Out & channel29_Kernel27_Valid_Out & channel30_Kernel27_Valid_Out & channel31_Kernel27_Valid_Out & channel32_Kernel27_Valid_Out & channel33_Kernel27_Valid_Out & channel34_Kernel27_Valid_Out & channel35_Kernel27_Valid_Out & channel36_Kernel27_Valid_Out & channel37_Kernel27_Valid_Out & channel38_Kernel27_Valid_Out & channel39_Kernel27_Valid_Out & channel40_Kernel27_Valid_Out & channel41_Kernel27_Valid_Out & channel42_Kernel27_Valid_Out & channel43_Kernel27_Valid_Out & channel44_Kernel27_Valid_Out & channel45_Kernel27_Valid_Out & channel46_Kernel27_Valid_Out & channel47_Kernel27_Valid_Out & channel48_Kernel27_Valid_Out & channel49_Kernel27_Valid_Out & channel50_Kernel27_Valid_Out & channel51_Kernel27_Valid_Out & channel52_Kernel27_Valid_Out & channel53_Kernel27_Valid_Out & channel54_Kernel27_Valid_Out & channel55_Kernel27_Valid_Out & channel56_Kernel27_Valid_Out & channel57_Kernel27_Valid_Out & channel58_Kernel27_Valid_Out & channel59_Kernel27_Valid_Out & channel60_Kernel27_Valid_Out & channel61_Kernel27_Valid_Out & channel62_Kernel27_Valid_Out & channel63_Kernel27_Valid_Out & channel64_Kernel27_Valid_Out;

	wire channel1_Kernel28_Valid_Out, channel2_Kernel28_Valid_Out, channel3_Kernel28_Valid_Out, channel4_Kernel28_Valid_Out, channel5_Kernel28_Valid_Out, channel6_Kernel28_Valid_Out, channel7_Kernel28_Valid_Out, channel8_Kernel28_Valid_Out, channel9_Kernel28_Valid_Out, channel10_Kernel28_Valid_Out, channel11_Kernel28_Valid_Out, channel12_Kernel28_Valid_Out, channel13_Kernel28_Valid_Out, channel14_Kernel28_Valid_Out, channel15_Kernel28_Valid_Out, channel16_Kernel28_Valid_Out, channel17_Kernel28_Valid_Out, channel18_Kernel28_Valid_Out, channel19_Kernel28_Valid_Out, channel20_Kernel28_Valid_Out, channel21_Kernel28_Valid_Out, channel22_Kernel28_Valid_Out, channel23_Kernel28_Valid_Out, channel24_Kernel28_Valid_Out, channel25_Kernel28_Valid_Out, channel26_Kernel28_Valid_Out, channel27_Kernel28_Valid_Out, channel28_Kernel28_Valid_Out, channel29_Kernel28_Valid_Out, channel30_Kernel28_Valid_Out, channel31_Kernel28_Valid_Out, channel32_Kernel28_Valid_Out, channel33_Kernel28_Valid_Out, channel34_Kernel28_Valid_Out, channel35_Kernel28_Valid_Out, channel36_Kernel28_Valid_Out, channel37_Kernel28_Valid_Out, channel38_Kernel28_Valid_Out, channel39_Kernel28_Valid_Out, channel40_Kernel28_Valid_Out, channel41_Kernel28_Valid_Out, channel42_Kernel28_Valid_Out, channel43_Kernel28_Valid_Out, channel44_Kernel28_Valid_Out, channel45_Kernel28_Valid_Out, channel46_Kernel28_Valid_Out, channel47_Kernel28_Valid_Out, channel48_Kernel28_Valid_Out, channel49_Kernel28_Valid_Out, channel50_Kernel28_Valid_Out, channel51_Kernel28_Valid_Out, channel52_Kernel28_Valid_Out, channel53_Kernel28_Valid_Out, channel54_Kernel28_Valid_Out, channel55_Kernel28_Valid_Out, channel56_Kernel28_Valid_Out, channel57_Kernel28_Valid_Out, channel58_Kernel28_Valid_Out, channel59_Kernel28_Valid_Out, channel60_Kernel28_Valid_Out, channel61_Kernel28_Valid_Out, channel62_Kernel28_Valid_Out, channel63_Kernel28_Valid_Out, channel64_Kernel28_Valid_Out;

	assign add_kernel28=channel1_Kernel28_Valid_Out & channel2_Kernel28_Valid_Out & channel3_Kernel28_Valid_Out & channel4_Kernel28_Valid_Out & channel5_Kernel28_Valid_Out & channel6_Kernel28_Valid_Out & channel7_Kernel28_Valid_Out & channel8_Kernel28_Valid_Out & channel9_Kernel28_Valid_Out & channel10_Kernel28_Valid_Out & channel11_Kernel28_Valid_Out & channel12_Kernel28_Valid_Out & channel13_Kernel28_Valid_Out & channel14_Kernel28_Valid_Out & channel15_Kernel28_Valid_Out & channel16_Kernel28_Valid_Out & channel17_Kernel28_Valid_Out & channel18_Kernel28_Valid_Out & channel19_Kernel28_Valid_Out & channel20_Kernel28_Valid_Out & channel21_Kernel28_Valid_Out & channel22_Kernel28_Valid_Out & channel23_Kernel28_Valid_Out & channel24_Kernel28_Valid_Out & channel25_Kernel28_Valid_Out & channel26_Kernel28_Valid_Out & channel27_Kernel28_Valid_Out & channel28_Kernel28_Valid_Out & channel29_Kernel28_Valid_Out & channel30_Kernel28_Valid_Out & channel31_Kernel28_Valid_Out & channel32_Kernel28_Valid_Out & channel33_Kernel28_Valid_Out & channel34_Kernel28_Valid_Out & channel35_Kernel28_Valid_Out & channel36_Kernel28_Valid_Out & channel37_Kernel28_Valid_Out & channel38_Kernel28_Valid_Out & channel39_Kernel28_Valid_Out & channel40_Kernel28_Valid_Out & channel41_Kernel28_Valid_Out & channel42_Kernel28_Valid_Out & channel43_Kernel28_Valid_Out & channel44_Kernel28_Valid_Out & channel45_Kernel28_Valid_Out & channel46_Kernel28_Valid_Out & channel47_Kernel28_Valid_Out & channel48_Kernel28_Valid_Out & channel49_Kernel28_Valid_Out & channel50_Kernel28_Valid_Out & channel51_Kernel28_Valid_Out & channel52_Kernel28_Valid_Out & channel53_Kernel28_Valid_Out & channel54_Kernel28_Valid_Out & channel55_Kernel28_Valid_Out & channel56_Kernel28_Valid_Out & channel57_Kernel28_Valid_Out & channel58_Kernel28_Valid_Out & channel59_Kernel28_Valid_Out & channel60_Kernel28_Valid_Out & channel61_Kernel28_Valid_Out & channel62_Kernel28_Valid_Out & channel63_Kernel28_Valid_Out & channel64_Kernel28_Valid_Out;

	wire channel1_Kernel29_Valid_Out, channel2_Kernel29_Valid_Out, channel3_Kernel29_Valid_Out, channel4_Kernel29_Valid_Out, channel5_Kernel29_Valid_Out, channel6_Kernel29_Valid_Out, channel7_Kernel29_Valid_Out, channel8_Kernel29_Valid_Out, channel9_Kernel29_Valid_Out, channel10_Kernel29_Valid_Out, channel11_Kernel29_Valid_Out, channel12_Kernel29_Valid_Out, channel13_Kernel29_Valid_Out, channel14_Kernel29_Valid_Out, channel15_Kernel29_Valid_Out, channel16_Kernel29_Valid_Out, channel17_Kernel29_Valid_Out, channel18_Kernel29_Valid_Out, channel19_Kernel29_Valid_Out, channel20_Kernel29_Valid_Out, channel21_Kernel29_Valid_Out, channel22_Kernel29_Valid_Out, channel23_Kernel29_Valid_Out, channel24_Kernel29_Valid_Out, channel25_Kernel29_Valid_Out, channel26_Kernel29_Valid_Out, channel27_Kernel29_Valid_Out, channel28_Kernel29_Valid_Out, channel29_Kernel29_Valid_Out, channel30_Kernel29_Valid_Out, channel31_Kernel29_Valid_Out, channel32_Kernel29_Valid_Out, channel33_Kernel29_Valid_Out, channel34_Kernel29_Valid_Out, channel35_Kernel29_Valid_Out, channel36_Kernel29_Valid_Out, channel37_Kernel29_Valid_Out, channel38_Kernel29_Valid_Out, channel39_Kernel29_Valid_Out, channel40_Kernel29_Valid_Out, channel41_Kernel29_Valid_Out, channel42_Kernel29_Valid_Out, channel43_Kernel29_Valid_Out, channel44_Kernel29_Valid_Out, channel45_Kernel29_Valid_Out, channel46_Kernel29_Valid_Out, channel47_Kernel29_Valid_Out, channel48_Kernel29_Valid_Out, channel49_Kernel29_Valid_Out, channel50_Kernel29_Valid_Out, channel51_Kernel29_Valid_Out, channel52_Kernel29_Valid_Out, channel53_Kernel29_Valid_Out, channel54_Kernel29_Valid_Out, channel55_Kernel29_Valid_Out, channel56_Kernel29_Valid_Out, channel57_Kernel29_Valid_Out, channel58_Kernel29_Valid_Out, channel59_Kernel29_Valid_Out, channel60_Kernel29_Valid_Out, channel61_Kernel29_Valid_Out, channel62_Kernel29_Valid_Out, channel63_Kernel29_Valid_Out, channel64_Kernel29_Valid_Out;

	assign add_kernel29=channel1_Kernel29_Valid_Out & channel2_Kernel29_Valid_Out & channel3_Kernel29_Valid_Out & channel4_Kernel29_Valid_Out & channel5_Kernel29_Valid_Out & channel6_Kernel29_Valid_Out & channel7_Kernel29_Valid_Out & channel8_Kernel29_Valid_Out & channel9_Kernel29_Valid_Out & channel10_Kernel29_Valid_Out & channel11_Kernel29_Valid_Out & channel12_Kernel29_Valid_Out & channel13_Kernel29_Valid_Out & channel14_Kernel29_Valid_Out & channel15_Kernel29_Valid_Out & channel16_Kernel29_Valid_Out & channel17_Kernel29_Valid_Out & channel18_Kernel29_Valid_Out & channel19_Kernel29_Valid_Out & channel20_Kernel29_Valid_Out & channel21_Kernel29_Valid_Out & channel22_Kernel29_Valid_Out & channel23_Kernel29_Valid_Out & channel24_Kernel29_Valid_Out & channel25_Kernel29_Valid_Out & channel26_Kernel29_Valid_Out & channel27_Kernel29_Valid_Out & channel28_Kernel29_Valid_Out & channel29_Kernel29_Valid_Out & channel30_Kernel29_Valid_Out & channel31_Kernel29_Valid_Out & channel32_Kernel29_Valid_Out & channel33_Kernel29_Valid_Out & channel34_Kernel29_Valid_Out & channel35_Kernel29_Valid_Out & channel36_Kernel29_Valid_Out & channel37_Kernel29_Valid_Out & channel38_Kernel29_Valid_Out & channel39_Kernel29_Valid_Out & channel40_Kernel29_Valid_Out & channel41_Kernel29_Valid_Out & channel42_Kernel29_Valid_Out & channel43_Kernel29_Valid_Out & channel44_Kernel29_Valid_Out & channel45_Kernel29_Valid_Out & channel46_Kernel29_Valid_Out & channel47_Kernel29_Valid_Out & channel48_Kernel29_Valid_Out & channel49_Kernel29_Valid_Out & channel50_Kernel29_Valid_Out & channel51_Kernel29_Valid_Out & channel52_Kernel29_Valid_Out & channel53_Kernel29_Valid_Out & channel54_Kernel29_Valid_Out & channel55_Kernel29_Valid_Out & channel56_Kernel29_Valid_Out & channel57_Kernel29_Valid_Out & channel58_Kernel29_Valid_Out & channel59_Kernel29_Valid_Out & channel60_Kernel29_Valid_Out & channel61_Kernel29_Valid_Out & channel62_Kernel29_Valid_Out & channel63_Kernel29_Valid_Out & channel64_Kernel29_Valid_Out;

	wire channel1_Kernel30_Valid_Out, channel2_Kernel30_Valid_Out, channel3_Kernel30_Valid_Out, channel4_Kernel30_Valid_Out, channel5_Kernel30_Valid_Out, channel6_Kernel30_Valid_Out, channel7_Kernel30_Valid_Out, channel8_Kernel30_Valid_Out, channel9_Kernel30_Valid_Out, channel10_Kernel30_Valid_Out, channel11_Kernel30_Valid_Out, channel12_Kernel30_Valid_Out, channel13_Kernel30_Valid_Out, channel14_Kernel30_Valid_Out, channel15_Kernel30_Valid_Out, channel16_Kernel30_Valid_Out, channel17_Kernel30_Valid_Out, channel18_Kernel30_Valid_Out, channel19_Kernel30_Valid_Out, channel20_Kernel30_Valid_Out, channel21_Kernel30_Valid_Out, channel22_Kernel30_Valid_Out, channel23_Kernel30_Valid_Out, channel24_Kernel30_Valid_Out, channel25_Kernel30_Valid_Out, channel26_Kernel30_Valid_Out, channel27_Kernel30_Valid_Out, channel28_Kernel30_Valid_Out, channel29_Kernel30_Valid_Out, channel30_Kernel30_Valid_Out, channel31_Kernel30_Valid_Out, channel32_Kernel30_Valid_Out, channel33_Kernel30_Valid_Out, channel34_Kernel30_Valid_Out, channel35_Kernel30_Valid_Out, channel36_Kernel30_Valid_Out, channel37_Kernel30_Valid_Out, channel38_Kernel30_Valid_Out, channel39_Kernel30_Valid_Out, channel40_Kernel30_Valid_Out, channel41_Kernel30_Valid_Out, channel42_Kernel30_Valid_Out, channel43_Kernel30_Valid_Out, channel44_Kernel30_Valid_Out, channel45_Kernel30_Valid_Out, channel46_Kernel30_Valid_Out, channel47_Kernel30_Valid_Out, channel48_Kernel30_Valid_Out, channel49_Kernel30_Valid_Out, channel50_Kernel30_Valid_Out, channel51_Kernel30_Valid_Out, channel52_Kernel30_Valid_Out, channel53_Kernel30_Valid_Out, channel54_Kernel30_Valid_Out, channel55_Kernel30_Valid_Out, channel56_Kernel30_Valid_Out, channel57_Kernel30_Valid_Out, channel58_Kernel30_Valid_Out, channel59_Kernel30_Valid_Out, channel60_Kernel30_Valid_Out, channel61_Kernel30_Valid_Out, channel62_Kernel30_Valid_Out, channel63_Kernel30_Valid_Out, channel64_Kernel30_Valid_Out;

	assign add_kernel30=channel1_Kernel30_Valid_Out & channel2_Kernel30_Valid_Out & channel3_Kernel30_Valid_Out & channel4_Kernel30_Valid_Out & channel5_Kernel30_Valid_Out & channel6_Kernel30_Valid_Out & channel7_Kernel30_Valid_Out & channel8_Kernel30_Valid_Out & channel9_Kernel30_Valid_Out & channel10_Kernel30_Valid_Out & channel11_Kernel30_Valid_Out & channel12_Kernel30_Valid_Out & channel13_Kernel30_Valid_Out & channel14_Kernel30_Valid_Out & channel15_Kernel30_Valid_Out & channel16_Kernel30_Valid_Out & channel17_Kernel30_Valid_Out & channel18_Kernel30_Valid_Out & channel19_Kernel30_Valid_Out & channel20_Kernel30_Valid_Out & channel21_Kernel30_Valid_Out & channel22_Kernel30_Valid_Out & channel23_Kernel30_Valid_Out & channel24_Kernel30_Valid_Out & channel25_Kernel30_Valid_Out & channel26_Kernel30_Valid_Out & channel27_Kernel30_Valid_Out & channel28_Kernel30_Valid_Out & channel29_Kernel30_Valid_Out & channel30_Kernel30_Valid_Out & channel31_Kernel30_Valid_Out & channel32_Kernel30_Valid_Out & channel33_Kernel30_Valid_Out & channel34_Kernel30_Valid_Out & channel35_Kernel30_Valid_Out & channel36_Kernel30_Valid_Out & channel37_Kernel30_Valid_Out & channel38_Kernel30_Valid_Out & channel39_Kernel30_Valid_Out & channel40_Kernel30_Valid_Out & channel41_Kernel30_Valid_Out & channel42_Kernel30_Valid_Out & channel43_Kernel30_Valid_Out & channel44_Kernel30_Valid_Out & channel45_Kernel30_Valid_Out & channel46_Kernel30_Valid_Out & channel47_Kernel30_Valid_Out & channel48_Kernel30_Valid_Out & channel49_Kernel30_Valid_Out & channel50_Kernel30_Valid_Out & channel51_Kernel30_Valid_Out & channel52_Kernel30_Valid_Out & channel53_Kernel30_Valid_Out & channel54_Kernel30_Valid_Out & channel55_Kernel30_Valid_Out & channel56_Kernel30_Valid_Out & channel57_Kernel30_Valid_Out & channel58_Kernel30_Valid_Out & channel59_Kernel30_Valid_Out & channel60_Kernel30_Valid_Out & channel61_Kernel30_Valid_Out & channel62_Kernel30_Valid_Out & channel63_Kernel30_Valid_Out & channel64_Kernel30_Valid_Out;

	wire channel1_Kernel31_Valid_Out, channel2_Kernel31_Valid_Out, channel3_Kernel31_Valid_Out, channel4_Kernel31_Valid_Out, channel5_Kernel31_Valid_Out, channel6_Kernel31_Valid_Out, channel7_Kernel31_Valid_Out, channel8_Kernel31_Valid_Out, channel9_Kernel31_Valid_Out, channel10_Kernel31_Valid_Out, channel11_Kernel31_Valid_Out, channel12_Kernel31_Valid_Out, channel13_Kernel31_Valid_Out, channel14_Kernel31_Valid_Out, channel15_Kernel31_Valid_Out, channel16_Kernel31_Valid_Out, channel17_Kernel31_Valid_Out, channel18_Kernel31_Valid_Out, channel19_Kernel31_Valid_Out, channel20_Kernel31_Valid_Out, channel21_Kernel31_Valid_Out, channel22_Kernel31_Valid_Out, channel23_Kernel31_Valid_Out, channel24_Kernel31_Valid_Out, channel25_Kernel31_Valid_Out, channel26_Kernel31_Valid_Out, channel27_Kernel31_Valid_Out, channel28_Kernel31_Valid_Out, channel29_Kernel31_Valid_Out, channel30_Kernel31_Valid_Out, channel31_Kernel31_Valid_Out, channel32_Kernel31_Valid_Out, channel33_Kernel31_Valid_Out, channel34_Kernel31_Valid_Out, channel35_Kernel31_Valid_Out, channel36_Kernel31_Valid_Out, channel37_Kernel31_Valid_Out, channel38_Kernel31_Valid_Out, channel39_Kernel31_Valid_Out, channel40_Kernel31_Valid_Out, channel41_Kernel31_Valid_Out, channel42_Kernel31_Valid_Out, channel43_Kernel31_Valid_Out, channel44_Kernel31_Valid_Out, channel45_Kernel31_Valid_Out, channel46_Kernel31_Valid_Out, channel47_Kernel31_Valid_Out, channel48_Kernel31_Valid_Out, channel49_Kernel31_Valid_Out, channel50_Kernel31_Valid_Out, channel51_Kernel31_Valid_Out, channel52_Kernel31_Valid_Out, channel53_Kernel31_Valid_Out, channel54_Kernel31_Valid_Out, channel55_Kernel31_Valid_Out, channel56_Kernel31_Valid_Out, channel57_Kernel31_Valid_Out, channel58_Kernel31_Valid_Out, channel59_Kernel31_Valid_Out, channel60_Kernel31_Valid_Out, channel61_Kernel31_Valid_Out, channel62_Kernel31_Valid_Out, channel63_Kernel31_Valid_Out, channel64_Kernel31_Valid_Out;

	assign add_kernel31=channel1_Kernel31_Valid_Out & channel2_Kernel31_Valid_Out & channel3_Kernel31_Valid_Out & channel4_Kernel31_Valid_Out & channel5_Kernel31_Valid_Out & channel6_Kernel31_Valid_Out & channel7_Kernel31_Valid_Out & channel8_Kernel31_Valid_Out & channel9_Kernel31_Valid_Out & channel10_Kernel31_Valid_Out & channel11_Kernel31_Valid_Out & channel12_Kernel31_Valid_Out & channel13_Kernel31_Valid_Out & channel14_Kernel31_Valid_Out & channel15_Kernel31_Valid_Out & channel16_Kernel31_Valid_Out & channel17_Kernel31_Valid_Out & channel18_Kernel31_Valid_Out & channel19_Kernel31_Valid_Out & channel20_Kernel31_Valid_Out & channel21_Kernel31_Valid_Out & channel22_Kernel31_Valid_Out & channel23_Kernel31_Valid_Out & channel24_Kernel31_Valid_Out & channel25_Kernel31_Valid_Out & channel26_Kernel31_Valid_Out & channel27_Kernel31_Valid_Out & channel28_Kernel31_Valid_Out & channel29_Kernel31_Valid_Out & channel30_Kernel31_Valid_Out & channel31_Kernel31_Valid_Out & channel32_Kernel31_Valid_Out & channel33_Kernel31_Valid_Out & channel34_Kernel31_Valid_Out & channel35_Kernel31_Valid_Out & channel36_Kernel31_Valid_Out & channel37_Kernel31_Valid_Out & channel38_Kernel31_Valid_Out & channel39_Kernel31_Valid_Out & channel40_Kernel31_Valid_Out & channel41_Kernel31_Valid_Out & channel42_Kernel31_Valid_Out & channel43_Kernel31_Valid_Out & channel44_Kernel31_Valid_Out & channel45_Kernel31_Valid_Out & channel46_Kernel31_Valid_Out & channel47_Kernel31_Valid_Out & channel48_Kernel31_Valid_Out & channel49_Kernel31_Valid_Out & channel50_Kernel31_Valid_Out & channel51_Kernel31_Valid_Out & channel52_Kernel31_Valid_Out & channel53_Kernel31_Valid_Out & channel54_Kernel31_Valid_Out & channel55_Kernel31_Valid_Out & channel56_Kernel31_Valid_Out & channel57_Kernel31_Valid_Out & channel58_Kernel31_Valid_Out & channel59_Kernel31_Valid_Out & channel60_Kernel31_Valid_Out & channel61_Kernel31_Valid_Out & channel62_Kernel31_Valid_Out & channel63_Kernel31_Valid_Out & channel64_Kernel31_Valid_Out;

	wire channel1_Kernel32_Valid_Out, channel2_Kernel32_Valid_Out, channel3_Kernel32_Valid_Out, channel4_Kernel32_Valid_Out, channel5_Kernel32_Valid_Out, channel6_Kernel32_Valid_Out, channel7_Kernel32_Valid_Out, channel8_Kernel32_Valid_Out, channel9_Kernel32_Valid_Out, channel10_Kernel32_Valid_Out, channel11_Kernel32_Valid_Out, channel12_Kernel32_Valid_Out, channel13_Kernel32_Valid_Out, channel14_Kernel32_Valid_Out, channel15_Kernel32_Valid_Out, channel16_Kernel32_Valid_Out, channel17_Kernel32_Valid_Out, channel18_Kernel32_Valid_Out, channel19_Kernel32_Valid_Out, channel20_Kernel32_Valid_Out, channel21_Kernel32_Valid_Out, channel22_Kernel32_Valid_Out, channel23_Kernel32_Valid_Out, channel24_Kernel32_Valid_Out, channel25_Kernel32_Valid_Out, channel26_Kernel32_Valid_Out, channel27_Kernel32_Valid_Out, channel28_Kernel32_Valid_Out, channel29_Kernel32_Valid_Out, channel30_Kernel32_Valid_Out, channel31_Kernel32_Valid_Out, channel32_Kernel32_Valid_Out, channel33_Kernel32_Valid_Out, channel34_Kernel32_Valid_Out, channel35_Kernel32_Valid_Out, channel36_Kernel32_Valid_Out, channel37_Kernel32_Valid_Out, channel38_Kernel32_Valid_Out, channel39_Kernel32_Valid_Out, channel40_Kernel32_Valid_Out, channel41_Kernel32_Valid_Out, channel42_Kernel32_Valid_Out, channel43_Kernel32_Valid_Out, channel44_Kernel32_Valid_Out, channel45_Kernel32_Valid_Out, channel46_Kernel32_Valid_Out, channel47_Kernel32_Valid_Out, channel48_Kernel32_Valid_Out, channel49_Kernel32_Valid_Out, channel50_Kernel32_Valid_Out, channel51_Kernel32_Valid_Out, channel52_Kernel32_Valid_Out, channel53_Kernel32_Valid_Out, channel54_Kernel32_Valid_Out, channel55_Kernel32_Valid_Out, channel56_Kernel32_Valid_Out, channel57_Kernel32_Valid_Out, channel58_Kernel32_Valid_Out, channel59_Kernel32_Valid_Out, channel60_Kernel32_Valid_Out, channel61_Kernel32_Valid_Out, channel62_Kernel32_Valid_Out, channel63_Kernel32_Valid_Out, channel64_Kernel32_Valid_Out;

	assign add_kernel32=channel1_Kernel32_Valid_Out & channel2_Kernel32_Valid_Out & channel3_Kernel32_Valid_Out & channel4_Kernel32_Valid_Out & channel5_Kernel32_Valid_Out & channel6_Kernel32_Valid_Out & channel7_Kernel32_Valid_Out & channel8_Kernel32_Valid_Out & channel9_Kernel32_Valid_Out & channel10_Kernel32_Valid_Out & channel11_Kernel32_Valid_Out & channel12_Kernel32_Valid_Out & channel13_Kernel32_Valid_Out & channel14_Kernel32_Valid_Out & channel15_Kernel32_Valid_Out & channel16_Kernel32_Valid_Out & channel17_Kernel32_Valid_Out & channel18_Kernel32_Valid_Out & channel19_Kernel32_Valid_Out & channel20_Kernel32_Valid_Out & channel21_Kernel32_Valid_Out & channel22_Kernel32_Valid_Out & channel23_Kernel32_Valid_Out & channel24_Kernel32_Valid_Out & channel25_Kernel32_Valid_Out & channel26_Kernel32_Valid_Out & channel27_Kernel32_Valid_Out & channel28_Kernel32_Valid_Out & channel29_Kernel32_Valid_Out & channel30_Kernel32_Valid_Out & channel31_Kernel32_Valid_Out & channel32_Kernel32_Valid_Out & channel33_Kernel32_Valid_Out & channel34_Kernel32_Valid_Out & channel35_Kernel32_Valid_Out & channel36_Kernel32_Valid_Out & channel37_Kernel32_Valid_Out & channel38_Kernel32_Valid_Out & channel39_Kernel32_Valid_Out & channel40_Kernel32_Valid_Out & channel41_Kernel32_Valid_Out & channel42_Kernel32_Valid_Out & channel43_Kernel32_Valid_Out & channel44_Kernel32_Valid_Out & channel45_Kernel32_Valid_Out & channel46_Kernel32_Valid_Out & channel47_Kernel32_Valid_Out & channel48_Kernel32_Valid_Out & channel49_Kernel32_Valid_Out & channel50_Kernel32_Valid_Out & channel51_Kernel32_Valid_Out & channel52_Kernel32_Valid_Out & channel53_Kernel32_Valid_Out & channel54_Kernel32_Valid_Out & channel55_Kernel32_Valid_Out & channel56_Kernel32_Valid_Out & channel57_Kernel32_Valid_Out & channel58_Kernel32_Valid_Out & channel59_Kernel32_Valid_Out & channel60_Kernel32_Valid_Out & channel61_Kernel32_Valid_Out & channel62_Kernel32_Valid_Out & channel63_Kernel32_Valid_Out & channel64_Kernel32_Valid_Out;

	wire channel1_Kernel33_Valid_Out, channel2_Kernel33_Valid_Out, channel3_Kernel33_Valid_Out, channel4_Kernel33_Valid_Out, channel5_Kernel33_Valid_Out, channel6_Kernel33_Valid_Out, channel7_Kernel33_Valid_Out, channel8_Kernel33_Valid_Out, channel9_Kernel33_Valid_Out, channel10_Kernel33_Valid_Out, channel11_Kernel33_Valid_Out, channel12_Kernel33_Valid_Out, channel13_Kernel33_Valid_Out, channel14_Kernel33_Valid_Out, channel15_Kernel33_Valid_Out, channel16_Kernel33_Valid_Out, channel17_Kernel33_Valid_Out, channel18_Kernel33_Valid_Out, channel19_Kernel33_Valid_Out, channel20_Kernel33_Valid_Out, channel21_Kernel33_Valid_Out, channel22_Kernel33_Valid_Out, channel23_Kernel33_Valid_Out, channel24_Kernel33_Valid_Out, channel25_Kernel33_Valid_Out, channel26_Kernel33_Valid_Out, channel27_Kernel33_Valid_Out, channel28_Kernel33_Valid_Out, channel29_Kernel33_Valid_Out, channel30_Kernel33_Valid_Out, channel31_Kernel33_Valid_Out, channel32_Kernel33_Valid_Out, channel33_Kernel33_Valid_Out, channel34_Kernel33_Valid_Out, channel35_Kernel33_Valid_Out, channel36_Kernel33_Valid_Out, channel37_Kernel33_Valid_Out, channel38_Kernel33_Valid_Out, channel39_Kernel33_Valid_Out, channel40_Kernel33_Valid_Out, channel41_Kernel33_Valid_Out, channel42_Kernel33_Valid_Out, channel43_Kernel33_Valid_Out, channel44_Kernel33_Valid_Out, channel45_Kernel33_Valid_Out, channel46_Kernel33_Valid_Out, channel47_Kernel33_Valid_Out, channel48_Kernel33_Valid_Out, channel49_Kernel33_Valid_Out, channel50_Kernel33_Valid_Out, channel51_Kernel33_Valid_Out, channel52_Kernel33_Valid_Out, channel53_Kernel33_Valid_Out, channel54_Kernel33_Valid_Out, channel55_Kernel33_Valid_Out, channel56_Kernel33_Valid_Out, channel57_Kernel33_Valid_Out, channel58_Kernel33_Valid_Out, channel59_Kernel33_Valid_Out, channel60_Kernel33_Valid_Out, channel61_Kernel33_Valid_Out, channel62_Kernel33_Valid_Out, channel63_Kernel33_Valid_Out, channel64_Kernel33_Valid_Out;

	assign add_kernel33=channel1_Kernel33_Valid_Out & channel2_Kernel33_Valid_Out & channel3_Kernel33_Valid_Out & channel4_Kernel33_Valid_Out & channel5_Kernel33_Valid_Out & channel6_Kernel33_Valid_Out & channel7_Kernel33_Valid_Out & channel8_Kernel33_Valid_Out & channel9_Kernel33_Valid_Out & channel10_Kernel33_Valid_Out & channel11_Kernel33_Valid_Out & channel12_Kernel33_Valid_Out & channel13_Kernel33_Valid_Out & channel14_Kernel33_Valid_Out & channel15_Kernel33_Valid_Out & channel16_Kernel33_Valid_Out & channel17_Kernel33_Valid_Out & channel18_Kernel33_Valid_Out & channel19_Kernel33_Valid_Out & channel20_Kernel33_Valid_Out & channel21_Kernel33_Valid_Out & channel22_Kernel33_Valid_Out & channel23_Kernel33_Valid_Out & channel24_Kernel33_Valid_Out & channel25_Kernel33_Valid_Out & channel26_Kernel33_Valid_Out & channel27_Kernel33_Valid_Out & channel28_Kernel33_Valid_Out & channel29_Kernel33_Valid_Out & channel30_Kernel33_Valid_Out & channel31_Kernel33_Valid_Out & channel32_Kernel33_Valid_Out & channel33_Kernel33_Valid_Out & channel34_Kernel33_Valid_Out & channel35_Kernel33_Valid_Out & channel36_Kernel33_Valid_Out & channel37_Kernel33_Valid_Out & channel38_Kernel33_Valid_Out & channel39_Kernel33_Valid_Out & channel40_Kernel33_Valid_Out & channel41_Kernel33_Valid_Out & channel42_Kernel33_Valid_Out & channel43_Kernel33_Valid_Out & channel44_Kernel33_Valid_Out & channel45_Kernel33_Valid_Out & channel46_Kernel33_Valid_Out & channel47_Kernel33_Valid_Out & channel48_Kernel33_Valid_Out & channel49_Kernel33_Valid_Out & channel50_Kernel33_Valid_Out & channel51_Kernel33_Valid_Out & channel52_Kernel33_Valid_Out & channel53_Kernel33_Valid_Out & channel54_Kernel33_Valid_Out & channel55_Kernel33_Valid_Out & channel56_Kernel33_Valid_Out & channel57_Kernel33_Valid_Out & channel58_Kernel33_Valid_Out & channel59_Kernel33_Valid_Out & channel60_Kernel33_Valid_Out & channel61_Kernel33_Valid_Out & channel62_Kernel33_Valid_Out & channel63_Kernel33_Valid_Out & channel64_Kernel33_Valid_Out;

	wire channel1_Kernel34_Valid_Out, channel2_Kernel34_Valid_Out, channel3_Kernel34_Valid_Out, channel4_Kernel34_Valid_Out, channel5_Kernel34_Valid_Out, channel6_Kernel34_Valid_Out, channel7_Kernel34_Valid_Out, channel8_Kernel34_Valid_Out, channel9_Kernel34_Valid_Out, channel10_Kernel34_Valid_Out, channel11_Kernel34_Valid_Out, channel12_Kernel34_Valid_Out, channel13_Kernel34_Valid_Out, channel14_Kernel34_Valid_Out, channel15_Kernel34_Valid_Out, channel16_Kernel34_Valid_Out, channel17_Kernel34_Valid_Out, channel18_Kernel34_Valid_Out, channel19_Kernel34_Valid_Out, channel20_Kernel34_Valid_Out, channel21_Kernel34_Valid_Out, channel22_Kernel34_Valid_Out, channel23_Kernel34_Valid_Out, channel24_Kernel34_Valid_Out, channel25_Kernel34_Valid_Out, channel26_Kernel34_Valid_Out, channel27_Kernel34_Valid_Out, channel28_Kernel34_Valid_Out, channel29_Kernel34_Valid_Out, channel30_Kernel34_Valid_Out, channel31_Kernel34_Valid_Out, channel32_Kernel34_Valid_Out, channel33_Kernel34_Valid_Out, channel34_Kernel34_Valid_Out, channel35_Kernel34_Valid_Out, channel36_Kernel34_Valid_Out, channel37_Kernel34_Valid_Out, channel38_Kernel34_Valid_Out, channel39_Kernel34_Valid_Out, channel40_Kernel34_Valid_Out, channel41_Kernel34_Valid_Out, channel42_Kernel34_Valid_Out, channel43_Kernel34_Valid_Out, channel44_Kernel34_Valid_Out, channel45_Kernel34_Valid_Out, channel46_Kernel34_Valid_Out, channel47_Kernel34_Valid_Out, channel48_Kernel34_Valid_Out, channel49_Kernel34_Valid_Out, channel50_Kernel34_Valid_Out, channel51_Kernel34_Valid_Out, channel52_Kernel34_Valid_Out, channel53_Kernel34_Valid_Out, channel54_Kernel34_Valid_Out, channel55_Kernel34_Valid_Out, channel56_Kernel34_Valid_Out, channel57_Kernel34_Valid_Out, channel58_Kernel34_Valid_Out, channel59_Kernel34_Valid_Out, channel60_Kernel34_Valid_Out, channel61_Kernel34_Valid_Out, channel62_Kernel34_Valid_Out, channel63_Kernel34_Valid_Out, channel64_Kernel34_Valid_Out;

	assign add_kernel34=channel1_Kernel34_Valid_Out & channel2_Kernel34_Valid_Out & channel3_Kernel34_Valid_Out & channel4_Kernel34_Valid_Out & channel5_Kernel34_Valid_Out & channel6_Kernel34_Valid_Out & channel7_Kernel34_Valid_Out & channel8_Kernel34_Valid_Out & channel9_Kernel34_Valid_Out & channel10_Kernel34_Valid_Out & channel11_Kernel34_Valid_Out & channel12_Kernel34_Valid_Out & channel13_Kernel34_Valid_Out & channel14_Kernel34_Valid_Out & channel15_Kernel34_Valid_Out & channel16_Kernel34_Valid_Out & channel17_Kernel34_Valid_Out & channel18_Kernel34_Valid_Out & channel19_Kernel34_Valid_Out & channel20_Kernel34_Valid_Out & channel21_Kernel34_Valid_Out & channel22_Kernel34_Valid_Out & channel23_Kernel34_Valid_Out & channel24_Kernel34_Valid_Out & channel25_Kernel34_Valid_Out & channel26_Kernel34_Valid_Out & channel27_Kernel34_Valid_Out & channel28_Kernel34_Valid_Out & channel29_Kernel34_Valid_Out & channel30_Kernel34_Valid_Out & channel31_Kernel34_Valid_Out & channel32_Kernel34_Valid_Out & channel33_Kernel34_Valid_Out & channel34_Kernel34_Valid_Out & channel35_Kernel34_Valid_Out & channel36_Kernel34_Valid_Out & channel37_Kernel34_Valid_Out & channel38_Kernel34_Valid_Out & channel39_Kernel34_Valid_Out & channel40_Kernel34_Valid_Out & channel41_Kernel34_Valid_Out & channel42_Kernel34_Valid_Out & channel43_Kernel34_Valid_Out & channel44_Kernel34_Valid_Out & channel45_Kernel34_Valid_Out & channel46_Kernel34_Valid_Out & channel47_Kernel34_Valid_Out & channel48_Kernel34_Valid_Out & channel49_Kernel34_Valid_Out & channel50_Kernel34_Valid_Out & channel51_Kernel34_Valid_Out & channel52_Kernel34_Valid_Out & channel53_Kernel34_Valid_Out & channel54_Kernel34_Valid_Out & channel55_Kernel34_Valid_Out & channel56_Kernel34_Valid_Out & channel57_Kernel34_Valid_Out & channel58_Kernel34_Valid_Out & channel59_Kernel34_Valid_Out & channel60_Kernel34_Valid_Out & channel61_Kernel34_Valid_Out & channel62_Kernel34_Valid_Out & channel63_Kernel34_Valid_Out & channel64_Kernel34_Valid_Out;

	wire channel1_Kernel35_Valid_Out, channel2_Kernel35_Valid_Out, channel3_Kernel35_Valid_Out, channel4_Kernel35_Valid_Out, channel5_Kernel35_Valid_Out, channel6_Kernel35_Valid_Out, channel7_Kernel35_Valid_Out, channel8_Kernel35_Valid_Out, channel9_Kernel35_Valid_Out, channel10_Kernel35_Valid_Out, channel11_Kernel35_Valid_Out, channel12_Kernel35_Valid_Out, channel13_Kernel35_Valid_Out, channel14_Kernel35_Valid_Out, channel15_Kernel35_Valid_Out, channel16_Kernel35_Valid_Out, channel17_Kernel35_Valid_Out, channel18_Kernel35_Valid_Out, channel19_Kernel35_Valid_Out, channel20_Kernel35_Valid_Out, channel21_Kernel35_Valid_Out, channel22_Kernel35_Valid_Out, channel23_Kernel35_Valid_Out, channel24_Kernel35_Valid_Out, channel25_Kernel35_Valid_Out, channel26_Kernel35_Valid_Out, channel27_Kernel35_Valid_Out, channel28_Kernel35_Valid_Out, channel29_Kernel35_Valid_Out, channel30_Kernel35_Valid_Out, channel31_Kernel35_Valid_Out, channel32_Kernel35_Valid_Out, channel33_Kernel35_Valid_Out, channel34_Kernel35_Valid_Out, channel35_Kernel35_Valid_Out, channel36_Kernel35_Valid_Out, channel37_Kernel35_Valid_Out, channel38_Kernel35_Valid_Out, channel39_Kernel35_Valid_Out, channel40_Kernel35_Valid_Out, channel41_Kernel35_Valid_Out, channel42_Kernel35_Valid_Out, channel43_Kernel35_Valid_Out, channel44_Kernel35_Valid_Out, channel45_Kernel35_Valid_Out, channel46_Kernel35_Valid_Out, channel47_Kernel35_Valid_Out, channel48_Kernel35_Valid_Out, channel49_Kernel35_Valid_Out, channel50_Kernel35_Valid_Out, channel51_Kernel35_Valid_Out, channel52_Kernel35_Valid_Out, channel53_Kernel35_Valid_Out, channel54_Kernel35_Valid_Out, channel55_Kernel35_Valid_Out, channel56_Kernel35_Valid_Out, channel57_Kernel35_Valid_Out, channel58_Kernel35_Valid_Out, channel59_Kernel35_Valid_Out, channel60_Kernel35_Valid_Out, channel61_Kernel35_Valid_Out, channel62_Kernel35_Valid_Out, channel63_Kernel35_Valid_Out, channel64_Kernel35_Valid_Out;

	assign add_kernel35=channel1_Kernel35_Valid_Out & channel2_Kernel35_Valid_Out & channel3_Kernel35_Valid_Out & channel4_Kernel35_Valid_Out & channel5_Kernel35_Valid_Out & channel6_Kernel35_Valid_Out & channel7_Kernel35_Valid_Out & channel8_Kernel35_Valid_Out & channel9_Kernel35_Valid_Out & channel10_Kernel35_Valid_Out & channel11_Kernel35_Valid_Out & channel12_Kernel35_Valid_Out & channel13_Kernel35_Valid_Out & channel14_Kernel35_Valid_Out & channel15_Kernel35_Valid_Out & channel16_Kernel35_Valid_Out & channel17_Kernel35_Valid_Out & channel18_Kernel35_Valid_Out & channel19_Kernel35_Valid_Out & channel20_Kernel35_Valid_Out & channel21_Kernel35_Valid_Out & channel22_Kernel35_Valid_Out & channel23_Kernel35_Valid_Out & channel24_Kernel35_Valid_Out & channel25_Kernel35_Valid_Out & channel26_Kernel35_Valid_Out & channel27_Kernel35_Valid_Out & channel28_Kernel35_Valid_Out & channel29_Kernel35_Valid_Out & channel30_Kernel35_Valid_Out & channel31_Kernel35_Valid_Out & channel32_Kernel35_Valid_Out & channel33_Kernel35_Valid_Out & channel34_Kernel35_Valid_Out & channel35_Kernel35_Valid_Out & channel36_Kernel35_Valid_Out & channel37_Kernel35_Valid_Out & channel38_Kernel35_Valid_Out & channel39_Kernel35_Valid_Out & channel40_Kernel35_Valid_Out & channel41_Kernel35_Valid_Out & channel42_Kernel35_Valid_Out & channel43_Kernel35_Valid_Out & channel44_Kernel35_Valid_Out & channel45_Kernel35_Valid_Out & channel46_Kernel35_Valid_Out & channel47_Kernel35_Valid_Out & channel48_Kernel35_Valid_Out & channel49_Kernel35_Valid_Out & channel50_Kernel35_Valid_Out & channel51_Kernel35_Valid_Out & channel52_Kernel35_Valid_Out & channel53_Kernel35_Valid_Out & channel54_Kernel35_Valid_Out & channel55_Kernel35_Valid_Out & channel56_Kernel35_Valid_Out & channel57_Kernel35_Valid_Out & channel58_Kernel35_Valid_Out & channel59_Kernel35_Valid_Out & channel60_Kernel35_Valid_Out & channel61_Kernel35_Valid_Out & channel62_Kernel35_Valid_Out & channel63_Kernel35_Valid_Out & channel64_Kernel35_Valid_Out;

	wire channel1_Kernel36_Valid_Out, channel2_Kernel36_Valid_Out, channel3_Kernel36_Valid_Out, channel4_Kernel36_Valid_Out, channel5_Kernel36_Valid_Out, channel6_Kernel36_Valid_Out, channel7_Kernel36_Valid_Out, channel8_Kernel36_Valid_Out, channel9_Kernel36_Valid_Out, channel10_Kernel36_Valid_Out, channel11_Kernel36_Valid_Out, channel12_Kernel36_Valid_Out, channel13_Kernel36_Valid_Out, channel14_Kernel36_Valid_Out, channel15_Kernel36_Valid_Out, channel16_Kernel36_Valid_Out, channel17_Kernel36_Valid_Out, channel18_Kernel36_Valid_Out, channel19_Kernel36_Valid_Out, channel20_Kernel36_Valid_Out, channel21_Kernel36_Valid_Out, channel22_Kernel36_Valid_Out, channel23_Kernel36_Valid_Out, channel24_Kernel36_Valid_Out, channel25_Kernel36_Valid_Out, channel26_Kernel36_Valid_Out, channel27_Kernel36_Valid_Out, channel28_Kernel36_Valid_Out, channel29_Kernel36_Valid_Out, channel30_Kernel36_Valid_Out, channel31_Kernel36_Valid_Out, channel32_Kernel36_Valid_Out, channel33_Kernel36_Valid_Out, channel34_Kernel36_Valid_Out, channel35_Kernel36_Valid_Out, channel36_Kernel36_Valid_Out, channel37_Kernel36_Valid_Out, channel38_Kernel36_Valid_Out, channel39_Kernel36_Valid_Out, channel40_Kernel36_Valid_Out, channel41_Kernel36_Valid_Out, channel42_Kernel36_Valid_Out, channel43_Kernel36_Valid_Out, channel44_Kernel36_Valid_Out, channel45_Kernel36_Valid_Out, channel46_Kernel36_Valid_Out, channel47_Kernel36_Valid_Out, channel48_Kernel36_Valid_Out, channel49_Kernel36_Valid_Out, channel50_Kernel36_Valid_Out, channel51_Kernel36_Valid_Out, channel52_Kernel36_Valid_Out, channel53_Kernel36_Valid_Out, channel54_Kernel36_Valid_Out, channel55_Kernel36_Valid_Out, channel56_Kernel36_Valid_Out, channel57_Kernel36_Valid_Out, channel58_Kernel36_Valid_Out, channel59_Kernel36_Valid_Out, channel60_Kernel36_Valid_Out, channel61_Kernel36_Valid_Out, channel62_Kernel36_Valid_Out, channel63_Kernel36_Valid_Out, channel64_Kernel36_Valid_Out;

	assign add_kernel36=channel1_Kernel36_Valid_Out & channel2_Kernel36_Valid_Out & channel3_Kernel36_Valid_Out & channel4_Kernel36_Valid_Out & channel5_Kernel36_Valid_Out & channel6_Kernel36_Valid_Out & channel7_Kernel36_Valid_Out & channel8_Kernel36_Valid_Out & channel9_Kernel36_Valid_Out & channel10_Kernel36_Valid_Out & channel11_Kernel36_Valid_Out & channel12_Kernel36_Valid_Out & channel13_Kernel36_Valid_Out & channel14_Kernel36_Valid_Out & channel15_Kernel36_Valid_Out & channel16_Kernel36_Valid_Out & channel17_Kernel36_Valid_Out & channel18_Kernel36_Valid_Out & channel19_Kernel36_Valid_Out & channel20_Kernel36_Valid_Out & channel21_Kernel36_Valid_Out & channel22_Kernel36_Valid_Out & channel23_Kernel36_Valid_Out & channel24_Kernel36_Valid_Out & channel25_Kernel36_Valid_Out & channel26_Kernel36_Valid_Out & channel27_Kernel36_Valid_Out & channel28_Kernel36_Valid_Out & channel29_Kernel36_Valid_Out & channel30_Kernel36_Valid_Out & channel31_Kernel36_Valid_Out & channel32_Kernel36_Valid_Out & channel33_Kernel36_Valid_Out & channel34_Kernel36_Valid_Out & channel35_Kernel36_Valid_Out & channel36_Kernel36_Valid_Out & channel37_Kernel36_Valid_Out & channel38_Kernel36_Valid_Out & channel39_Kernel36_Valid_Out & channel40_Kernel36_Valid_Out & channel41_Kernel36_Valid_Out & channel42_Kernel36_Valid_Out & channel43_Kernel36_Valid_Out & channel44_Kernel36_Valid_Out & channel45_Kernel36_Valid_Out & channel46_Kernel36_Valid_Out & channel47_Kernel36_Valid_Out & channel48_Kernel36_Valid_Out & channel49_Kernel36_Valid_Out & channel50_Kernel36_Valid_Out & channel51_Kernel36_Valid_Out & channel52_Kernel36_Valid_Out & channel53_Kernel36_Valid_Out & channel54_Kernel36_Valid_Out & channel55_Kernel36_Valid_Out & channel56_Kernel36_Valid_Out & channel57_Kernel36_Valid_Out & channel58_Kernel36_Valid_Out & channel59_Kernel36_Valid_Out & channel60_Kernel36_Valid_Out & channel61_Kernel36_Valid_Out & channel62_Kernel36_Valid_Out & channel63_Kernel36_Valid_Out & channel64_Kernel36_Valid_Out;

	wire channel1_Kernel37_Valid_Out, channel2_Kernel37_Valid_Out, channel3_Kernel37_Valid_Out, channel4_Kernel37_Valid_Out, channel5_Kernel37_Valid_Out, channel6_Kernel37_Valid_Out, channel7_Kernel37_Valid_Out, channel8_Kernel37_Valid_Out, channel9_Kernel37_Valid_Out, channel10_Kernel37_Valid_Out, channel11_Kernel37_Valid_Out, channel12_Kernel37_Valid_Out, channel13_Kernel37_Valid_Out, channel14_Kernel37_Valid_Out, channel15_Kernel37_Valid_Out, channel16_Kernel37_Valid_Out, channel17_Kernel37_Valid_Out, channel18_Kernel37_Valid_Out, channel19_Kernel37_Valid_Out, channel20_Kernel37_Valid_Out, channel21_Kernel37_Valid_Out, channel22_Kernel37_Valid_Out, channel23_Kernel37_Valid_Out, channel24_Kernel37_Valid_Out, channel25_Kernel37_Valid_Out, channel26_Kernel37_Valid_Out, channel27_Kernel37_Valid_Out, channel28_Kernel37_Valid_Out, channel29_Kernel37_Valid_Out, channel30_Kernel37_Valid_Out, channel31_Kernel37_Valid_Out, channel32_Kernel37_Valid_Out, channel33_Kernel37_Valid_Out, channel34_Kernel37_Valid_Out, channel35_Kernel37_Valid_Out, channel36_Kernel37_Valid_Out, channel37_Kernel37_Valid_Out, channel38_Kernel37_Valid_Out, channel39_Kernel37_Valid_Out, channel40_Kernel37_Valid_Out, channel41_Kernel37_Valid_Out, channel42_Kernel37_Valid_Out, channel43_Kernel37_Valid_Out, channel44_Kernel37_Valid_Out, channel45_Kernel37_Valid_Out, channel46_Kernel37_Valid_Out, channel47_Kernel37_Valid_Out, channel48_Kernel37_Valid_Out, channel49_Kernel37_Valid_Out, channel50_Kernel37_Valid_Out, channel51_Kernel37_Valid_Out, channel52_Kernel37_Valid_Out, channel53_Kernel37_Valid_Out, channel54_Kernel37_Valid_Out, channel55_Kernel37_Valid_Out, channel56_Kernel37_Valid_Out, channel57_Kernel37_Valid_Out, channel58_Kernel37_Valid_Out, channel59_Kernel37_Valid_Out, channel60_Kernel37_Valid_Out, channel61_Kernel37_Valid_Out, channel62_Kernel37_Valid_Out, channel63_Kernel37_Valid_Out, channel64_Kernel37_Valid_Out;

	assign add_kernel37=channel1_Kernel37_Valid_Out & channel2_Kernel37_Valid_Out & channel3_Kernel37_Valid_Out & channel4_Kernel37_Valid_Out & channel5_Kernel37_Valid_Out & channel6_Kernel37_Valid_Out & channel7_Kernel37_Valid_Out & channel8_Kernel37_Valid_Out & channel9_Kernel37_Valid_Out & channel10_Kernel37_Valid_Out & channel11_Kernel37_Valid_Out & channel12_Kernel37_Valid_Out & channel13_Kernel37_Valid_Out & channel14_Kernel37_Valid_Out & channel15_Kernel37_Valid_Out & channel16_Kernel37_Valid_Out & channel17_Kernel37_Valid_Out & channel18_Kernel37_Valid_Out & channel19_Kernel37_Valid_Out & channel20_Kernel37_Valid_Out & channel21_Kernel37_Valid_Out & channel22_Kernel37_Valid_Out & channel23_Kernel37_Valid_Out & channel24_Kernel37_Valid_Out & channel25_Kernel37_Valid_Out & channel26_Kernel37_Valid_Out & channel27_Kernel37_Valid_Out & channel28_Kernel37_Valid_Out & channel29_Kernel37_Valid_Out & channel30_Kernel37_Valid_Out & channel31_Kernel37_Valid_Out & channel32_Kernel37_Valid_Out & channel33_Kernel37_Valid_Out & channel34_Kernel37_Valid_Out & channel35_Kernel37_Valid_Out & channel36_Kernel37_Valid_Out & channel37_Kernel37_Valid_Out & channel38_Kernel37_Valid_Out & channel39_Kernel37_Valid_Out & channel40_Kernel37_Valid_Out & channel41_Kernel37_Valid_Out & channel42_Kernel37_Valid_Out & channel43_Kernel37_Valid_Out & channel44_Kernel37_Valid_Out & channel45_Kernel37_Valid_Out & channel46_Kernel37_Valid_Out & channel47_Kernel37_Valid_Out & channel48_Kernel37_Valid_Out & channel49_Kernel37_Valid_Out & channel50_Kernel37_Valid_Out & channel51_Kernel37_Valid_Out & channel52_Kernel37_Valid_Out & channel53_Kernel37_Valid_Out & channel54_Kernel37_Valid_Out & channel55_Kernel37_Valid_Out & channel56_Kernel37_Valid_Out & channel57_Kernel37_Valid_Out & channel58_Kernel37_Valid_Out & channel59_Kernel37_Valid_Out & channel60_Kernel37_Valid_Out & channel61_Kernel37_Valid_Out & channel62_Kernel37_Valid_Out & channel63_Kernel37_Valid_Out & channel64_Kernel37_Valid_Out;

	wire channel1_Kernel38_Valid_Out, channel2_Kernel38_Valid_Out, channel3_Kernel38_Valid_Out, channel4_Kernel38_Valid_Out, channel5_Kernel38_Valid_Out, channel6_Kernel38_Valid_Out, channel7_Kernel38_Valid_Out, channel8_Kernel38_Valid_Out, channel9_Kernel38_Valid_Out, channel10_Kernel38_Valid_Out, channel11_Kernel38_Valid_Out, channel12_Kernel38_Valid_Out, channel13_Kernel38_Valid_Out, channel14_Kernel38_Valid_Out, channel15_Kernel38_Valid_Out, channel16_Kernel38_Valid_Out, channel17_Kernel38_Valid_Out, channel18_Kernel38_Valid_Out, channel19_Kernel38_Valid_Out, channel20_Kernel38_Valid_Out, channel21_Kernel38_Valid_Out, channel22_Kernel38_Valid_Out, channel23_Kernel38_Valid_Out, channel24_Kernel38_Valid_Out, channel25_Kernel38_Valid_Out, channel26_Kernel38_Valid_Out, channel27_Kernel38_Valid_Out, channel28_Kernel38_Valid_Out, channel29_Kernel38_Valid_Out, channel30_Kernel38_Valid_Out, channel31_Kernel38_Valid_Out, channel32_Kernel38_Valid_Out, channel33_Kernel38_Valid_Out, channel34_Kernel38_Valid_Out, channel35_Kernel38_Valid_Out, channel36_Kernel38_Valid_Out, channel37_Kernel38_Valid_Out, channel38_Kernel38_Valid_Out, channel39_Kernel38_Valid_Out, channel40_Kernel38_Valid_Out, channel41_Kernel38_Valid_Out, channel42_Kernel38_Valid_Out, channel43_Kernel38_Valid_Out, channel44_Kernel38_Valid_Out, channel45_Kernel38_Valid_Out, channel46_Kernel38_Valid_Out, channel47_Kernel38_Valid_Out, channel48_Kernel38_Valid_Out, channel49_Kernel38_Valid_Out, channel50_Kernel38_Valid_Out, channel51_Kernel38_Valid_Out, channel52_Kernel38_Valid_Out, channel53_Kernel38_Valid_Out, channel54_Kernel38_Valid_Out, channel55_Kernel38_Valid_Out, channel56_Kernel38_Valid_Out, channel57_Kernel38_Valid_Out, channel58_Kernel38_Valid_Out, channel59_Kernel38_Valid_Out, channel60_Kernel38_Valid_Out, channel61_Kernel38_Valid_Out, channel62_Kernel38_Valid_Out, channel63_Kernel38_Valid_Out, channel64_Kernel38_Valid_Out;

	assign add_kernel38=channel1_Kernel38_Valid_Out & channel2_Kernel38_Valid_Out & channel3_Kernel38_Valid_Out & channel4_Kernel38_Valid_Out & channel5_Kernel38_Valid_Out & channel6_Kernel38_Valid_Out & channel7_Kernel38_Valid_Out & channel8_Kernel38_Valid_Out & channel9_Kernel38_Valid_Out & channel10_Kernel38_Valid_Out & channel11_Kernel38_Valid_Out & channel12_Kernel38_Valid_Out & channel13_Kernel38_Valid_Out & channel14_Kernel38_Valid_Out & channel15_Kernel38_Valid_Out & channel16_Kernel38_Valid_Out & channel17_Kernel38_Valid_Out & channel18_Kernel38_Valid_Out & channel19_Kernel38_Valid_Out & channel20_Kernel38_Valid_Out & channel21_Kernel38_Valid_Out & channel22_Kernel38_Valid_Out & channel23_Kernel38_Valid_Out & channel24_Kernel38_Valid_Out & channel25_Kernel38_Valid_Out & channel26_Kernel38_Valid_Out & channel27_Kernel38_Valid_Out & channel28_Kernel38_Valid_Out & channel29_Kernel38_Valid_Out & channel30_Kernel38_Valid_Out & channel31_Kernel38_Valid_Out & channel32_Kernel38_Valid_Out & channel33_Kernel38_Valid_Out & channel34_Kernel38_Valid_Out & channel35_Kernel38_Valid_Out & channel36_Kernel38_Valid_Out & channel37_Kernel38_Valid_Out & channel38_Kernel38_Valid_Out & channel39_Kernel38_Valid_Out & channel40_Kernel38_Valid_Out & channel41_Kernel38_Valid_Out & channel42_Kernel38_Valid_Out & channel43_Kernel38_Valid_Out & channel44_Kernel38_Valid_Out & channel45_Kernel38_Valid_Out & channel46_Kernel38_Valid_Out & channel47_Kernel38_Valid_Out & channel48_Kernel38_Valid_Out & channel49_Kernel38_Valid_Out & channel50_Kernel38_Valid_Out & channel51_Kernel38_Valid_Out & channel52_Kernel38_Valid_Out & channel53_Kernel38_Valid_Out & channel54_Kernel38_Valid_Out & channel55_Kernel38_Valid_Out & channel56_Kernel38_Valid_Out & channel57_Kernel38_Valid_Out & channel58_Kernel38_Valid_Out & channel59_Kernel38_Valid_Out & channel60_Kernel38_Valid_Out & channel61_Kernel38_Valid_Out & channel62_Kernel38_Valid_Out & channel63_Kernel38_Valid_Out & channel64_Kernel38_Valid_Out;

	wire channel1_Kernel39_Valid_Out, channel2_Kernel39_Valid_Out, channel3_Kernel39_Valid_Out, channel4_Kernel39_Valid_Out, channel5_Kernel39_Valid_Out, channel6_Kernel39_Valid_Out, channel7_Kernel39_Valid_Out, channel8_Kernel39_Valid_Out, channel9_Kernel39_Valid_Out, channel10_Kernel39_Valid_Out, channel11_Kernel39_Valid_Out, channel12_Kernel39_Valid_Out, channel13_Kernel39_Valid_Out, channel14_Kernel39_Valid_Out, channel15_Kernel39_Valid_Out, channel16_Kernel39_Valid_Out, channel17_Kernel39_Valid_Out, channel18_Kernel39_Valid_Out, channel19_Kernel39_Valid_Out, channel20_Kernel39_Valid_Out, channel21_Kernel39_Valid_Out, channel22_Kernel39_Valid_Out, channel23_Kernel39_Valid_Out, channel24_Kernel39_Valid_Out, channel25_Kernel39_Valid_Out, channel26_Kernel39_Valid_Out, channel27_Kernel39_Valid_Out, channel28_Kernel39_Valid_Out, channel29_Kernel39_Valid_Out, channel30_Kernel39_Valid_Out, channel31_Kernel39_Valid_Out, channel32_Kernel39_Valid_Out, channel33_Kernel39_Valid_Out, channel34_Kernel39_Valid_Out, channel35_Kernel39_Valid_Out, channel36_Kernel39_Valid_Out, channel37_Kernel39_Valid_Out, channel38_Kernel39_Valid_Out, channel39_Kernel39_Valid_Out, channel40_Kernel39_Valid_Out, channel41_Kernel39_Valid_Out, channel42_Kernel39_Valid_Out, channel43_Kernel39_Valid_Out, channel44_Kernel39_Valid_Out, channel45_Kernel39_Valid_Out, channel46_Kernel39_Valid_Out, channel47_Kernel39_Valid_Out, channel48_Kernel39_Valid_Out, channel49_Kernel39_Valid_Out, channel50_Kernel39_Valid_Out, channel51_Kernel39_Valid_Out, channel52_Kernel39_Valid_Out, channel53_Kernel39_Valid_Out, channel54_Kernel39_Valid_Out, channel55_Kernel39_Valid_Out, channel56_Kernel39_Valid_Out, channel57_Kernel39_Valid_Out, channel58_Kernel39_Valid_Out, channel59_Kernel39_Valid_Out, channel60_Kernel39_Valid_Out, channel61_Kernel39_Valid_Out, channel62_Kernel39_Valid_Out, channel63_Kernel39_Valid_Out, channel64_Kernel39_Valid_Out;

	assign add_kernel39=channel1_Kernel39_Valid_Out & channel2_Kernel39_Valid_Out & channel3_Kernel39_Valid_Out & channel4_Kernel39_Valid_Out & channel5_Kernel39_Valid_Out & channel6_Kernel39_Valid_Out & channel7_Kernel39_Valid_Out & channel8_Kernel39_Valid_Out & channel9_Kernel39_Valid_Out & channel10_Kernel39_Valid_Out & channel11_Kernel39_Valid_Out & channel12_Kernel39_Valid_Out & channel13_Kernel39_Valid_Out & channel14_Kernel39_Valid_Out & channel15_Kernel39_Valid_Out & channel16_Kernel39_Valid_Out & channel17_Kernel39_Valid_Out & channel18_Kernel39_Valid_Out & channel19_Kernel39_Valid_Out & channel20_Kernel39_Valid_Out & channel21_Kernel39_Valid_Out & channel22_Kernel39_Valid_Out & channel23_Kernel39_Valid_Out & channel24_Kernel39_Valid_Out & channel25_Kernel39_Valid_Out & channel26_Kernel39_Valid_Out & channel27_Kernel39_Valid_Out & channel28_Kernel39_Valid_Out & channel29_Kernel39_Valid_Out & channel30_Kernel39_Valid_Out & channel31_Kernel39_Valid_Out & channel32_Kernel39_Valid_Out & channel33_Kernel39_Valid_Out & channel34_Kernel39_Valid_Out & channel35_Kernel39_Valid_Out & channel36_Kernel39_Valid_Out & channel37_Kernel39_Valid_Out & channel38_Kernel39_Valid_Out & channel39_Kernel39_Valid_Out & channel40_Kernel39_Valid_Out & channel41_Kernel39_Valid_Out & channel42_Kernel39_Valid_Out & channel43_Kernel39_Valid_Out & channel44_Kernel39_Valid_Out & channel45_Kernel39_Valid_Out & channel46_Kernel39_Valid_Out & channel47_Kernel39_Valid_Out & channel48_Kernel39_Valid_Out & channel49_Kernel39_Valid_Out & channel50_Kernel39_Valid_Out & channel51_Kernel39_Valid_Out & channel52_Kernel39_Valid_Out & channel53_Kernel39_Valid_Out & channel54_Kernel39_Valid_Out & channel55_Kernel39_Valid_Out & channel56_Kernel39_Valid_Out & channel57_Kernel39_Valid_Out & channel58_Kernel39_Valid_Out & channel59_Kernel39_Valid_Out & channel60_Kernel39_Valid_Out & channel61_Kernel39_Valid_Out & channel62_Kernel39_Valid_Out & channel63_Kernel39_Valid_Out & channel64_Kernel39_Valid_Out;

	wire channel1_Kernel40_Valid_Out, channel2_Kernel40_Valid_Out, channel3_Kernel40_Valid_Out, channel4_Kernel40_Valid_Out, channel5_Kernel40_Valid_Out, channel6_Kernel40_Valid_Out, channel7_Kernel40_Valid_Out, channel8_Kernel40_Valid_Out, channel9_Kernel40_Valid_Out, channel10_Kernel40_Valid_Out, channel11_Kernel40_Valid_Out, channel12_Kernel40_Valid_Out, channel13_Kernel40_Valid_Out, channel14_Kernel40_Valid_Out, channel15_Kernel40_Valid_Out, channel16_Kernel40_Valid_Out, channel17_Kernel40_Valid_Out, channel18_Kernel40_Valid_Out, channel19_Kernel40_Valid_Out, channel20_Kernel40_Valid_Out, channel21_Kernel40_Valid_Out, channel22_Kernel40_Valid_Out, channel23_Kernel40_Valid_Out, channel24_Kernel40_Valid_Out, channel25_Kernel40_Valid_Out, channel26_Kernel40_Valid_Out, channel27_Kernel40_Valid_Out, channel28_Kernel40_Valid_Out, channel29_Kernel40_Valid_Out, channel30_Kernel40_Valid_Out, channel31_Kernel40_Valid_Out, channel32_Kernel40_Valid_Out, channel33_Kernel40_Valid_Out, channel34_Kernel40_Valid_Out, channel35_Kernel40_Valid_Out, channel36_Kernel40_Valid_Out, channel37_Kernel40_Valid_Out, channel38_Kernel40_Valid_Out, channel39_Kernel40_Valid_Out, channel40_Kernel40_Valid_Out, channel41_Kernel40_Valid_Out, channel42_Kernel40_Valid_Out, channel43_Kernel40_Valid_Out, channel44_Kernel40_Valid_Out, channel45_Kernel40_Valid_Out, channel46_Kernel40_Valid_Out, channel47_Kernel40_Valid_Out, channel48_Kernel40_Valid_Out, channel49_Kernel40_Valid_Out, channel50_Kernel40_Valid_Out, channel51_Kernel40_Valid_Out, channel52_Kernel40_Valid_Out, channel53_Kernel40_Valid_Out, channel54_Kernel40_Valid_Out, channel55_Kernel40_Valid_Out, channel56_Kernel40_Valid_Out, channel57_Kernel40_Valid_Out, channel58_Kernel40_Valid_Out, channel59_Kernel40_Valid_Out, channel60_Kernel40_Valid_Out, channel61_Kernel40_Valid_Out, channel62_Kernel40_Valid_Out, channel63_Kernel40_Valid_Out, channel64_Kernel40_Valid_Out;

	assign add_kernel40=channel1_Kernel40_Valid_Out & channel2_Kernel40_Valid_Out & channel3_Kernel40_Valid_Out & channel4_Kernel40_Valid_Out & channel5_Kernel40_Valid_Out & channel6_Kernel40_Valid_Out & channel7_Kernel40_Valid_Out & channel8_Kernel40_Valid_Out & channel9_Kernel40_Valid_Out & channel10_Kernel40_Valid_Out & channel11_Kernel40_Valid_Out & channel12_Kernel40_Valid_Out & channel13_Kernel40_Valid_Out & channel14_Kernel40_Valid_Out & channel15_Kernel40_Valid_Out & channel16_Kernel40_Valid_Out & channel17_Kernel40_Valid_Out & channel18_Kernel40_Valid_Out & channel19_Kernel40_Valid_Out & channel20_Kernel40_Valid_Out & channel21_Kernel40_Valid_Out & channel22_Kernel40_Valid_Out & channel23_Kernel40_Valid_Out & channel24_Kernel40_Valid_Out & channel25_Kernel40_Valid_Out & channel26_Kernel40_Valid_Out & channel27_Kernel40_Valid_Out & channel28_Kernel40_Valid_Out & channel29_Kernel40_Valid_Out & channel30_Kernel40_Valid_Out & channel31_Kernel40_Valid_Out & channel32_Kernel40_Valid_Out & channel33_Kernel40_Valid_Out & channel34_Kernel40_Valid_Out & channel35_Kernel40_Valid_Out & channel36_Kernel40_Valid_Out & channel37_Kernel40_Valid_Out & channel38_Kernel40_Valid_Out & channel39_Kernel40_Valid_Out & channel40_Kernel40_Valid_Out & channel41_Kernel40_Valid_Out & channel42_Kernel40_Valid_Out & channel43_Kernel40_Valid_Out & channel44_Kernel40_Valid_Out & channel45_Kernel40_Valid_Out & channel46_Kernel40_Valid_Out & channel47_Kernel40_Valid_Out & channel48_Kernel40_Valid_Out & channel49_Kernel40_Valid_Out & channel50_Kernel40_Valid_Out & channel51_Kernel40_Valid_Out & channel52_Kernel40_Valid_Out & channel53_Kernel40_Valid_Out & channel54_Kernel40_Valid_Out & channel55_Kernel40_Valid_Out & channel56_Kernel40_Valid_Out & channel57_Kernel40_Valid_Out & channel58_Kernel40_Valid_Out & channel59_Kernel40_Valid_Out & channel60_Kernel40_Valid_Out & channel61_Kernel40_Valid_Out & channel62_Kernel40_Valid_Out & channel63_Kernel40_Valid_Out & channel64_Kernel40_Valid_Out;

	wire channel1_Kernel41_Valid_Out, channel2_Kernel41_Valid_Out, channel3_Kernel41_Valid_Out, channel4_Kernel41_Valid_Out, channel5_Kernel41_Valid_Out, channel6_Kernel41_Valid_Out, channel7_Kernel41_Valid_Out, channel8_Kernel41_Valid_Out, channel9_Kernel41_Valid_Out, channel10_Kernel41_Valid_Out, channel11_Kernel41_Valid_Out, channel12_Kernel41_Valid_Out, channel13_Kernel41_Valid_Out, channel14_Kernel41_Valid_Out, channel15_Kernel41_Valid_Out, channel16_Kernel41_Valid_Out, channel17_Kernel41_Valid_Out, channel18_Kernel41_Valid_Out, channel19_Kernel41_Valid_Out, channel20_Kernel41_Valid_Out, channel21_Kernel41_Valid_Out, channel22_Kernel41_Valid_Out, channel23_Kernel41_Valid_Out, channel24_Kernel41_Valid_Out, channel25_Kernel41_Valid_Out, channel26_Kernel41_Valid_Out, channel27_Kernel41_Valid_Out, channel28_Kernel41_Valid_Out, channel29_Kernel41_Valid_Out, channel30_Kernel41_Valid_Out, channel31_Kernel41_Valid_Out, channel32_Kernel41_Valid_Out, channel33_Kernel41_Valid_Out, channel34_Kernel41_Valid_Out, channel35_Kernel41_Valid_Out, channel36_Kernel41_Valid_Out, channel37_Kernel41_Valid_Out, channel38_Kernel41_Valid_Out, channel39_Kernel41_Valid_Out, channel40_Kernel41_Valid_Out, channel41_Kernel41_Valid_Out, channel42_Kernel41_Valid_Out, channel43_Kernel41_Valid_Out, channel44_Kernel41_Valid_Out, channel45_Kernel41_Valid_Out, channel46_Kernel41_Valid_Out, channel47_Kernel41_Valid_Out, channel48_Kernel41_Valid_Out, channel49_Kernel41_Valid_Out, channel50_Kernel41_Valid_Out, channel51_Kernel41_Valid_Out, channel52_Kernel41_Valid_Out, channel53_Kernel41_Valid_Out, channel54_Kernel41_Valid_Out, channel55_Kernel41_Valid_Out, channel56_Kernel41_Valid_Out, channel57_Kernel41_Valid_Out, channel58_Kernel41_Valid_Out, channel59_Kernel41_Valid_Out, channel60_Kernel41_Valid_Out, channel61_Kernel41_Valid_Out, channel62_Kernel41_Valid_Out, channel63_Kernel41_Valid_Out, channel64_Kernel41_Valid_Out;

	assign add_kernel41=channel1_Kernel41_Valid_Out & channel2_Kernel41_Valid_Out & channel3_Kernel41_Valid_Out & channel4_Kernel41_Valid_Out & channel5_Kernel41_Valid_Out & channel6_Kernel41_Valid_Out & channel7_Kernel41_Valid_Out & channel8_Kernel41_Valid_Out & channel9_Kernel41_Valid_Out & channel10_Kernel41_Valid_Out & channel11_Kernel41_Valid_Out & channel12_Kernel41_Valid_Out & channel13_Kernel41_Valid_Out & channel14_Kernel41_Valid_Out & channel15_Kernel41_Valid_Out & channel16_Kernel41_Valid_Out & channel17_Kernel41_Valid_Out & channel18_Kernel41_Valid_Out & channel19_Kernel41_Valid_Out & channel20_Kernel41_Valid_Out & channel21_Kernel41_Valid_Out & channel22_Kernel41_Valid_Out & channel23_Kernel41_Valid_Out & channel24_Kernel41_Valid_Out & channel25_Kernel41_Valid_Out & channel26_Kernel41_Valid_Out & channel27_Kernel41_Valid_Out & channel28_Kernel41_Valid_Out & channel29_Kernel41_Valid_Out & channel30_Kernel41_Valid_Out & channel31_Kernel41_Valid_Out & channel32_Kernel41_Valid_Out & channel33_Kernel41_Valid_Out & channel34_Kernel41_Valid_Out & channel35_Kernel41_Valid_Out & channel36_Kernel41_Valid_Out & channel37_Kernel41_Valid_Out & channel38_Kernel41_Valid_Out & channel39_Kernel41_Valid_Out & channel40_Kernel41_Valid_Out & channel41_Kernel41_Valid_Out & channel42_Kernel41_Valid_Out & channel43_Kernel41_Valid_Out & channel44_Kernel41_Valid_Out & channel45_Kernel41_Valid_Out & channel46_Kernel41_Valid_Out & channel47_Kernel41_Valid_Out & channel48_Kernel41_Valid_Out & channel49_Kernel41_Valid_Out & channel50_Kernel41_Valid_Out & channel51_Kernel41_Valid_Out & channel52_Kernel41_Valid_Out & channel53_Kernel41_Valid_Out & channel54_Kernel41_Valid_Out & channel55_Kernel41_Valid_Out & channel56_Kernel41_Valid_Out & channel57_Kernel41_Valid_Out & channel58_Kernel41_Valid_Out & channel59_Kernel41_Valid_Out & channel60_Kernel41_Valid_Out & channel61_Kernel41_Valid_Out & channel62_Kernel41_Valid_Out & channel63_Kernel41_Valid_Out & channel64_Kernel41_Valid_Out;

	wire channel1_Kernel42_Valid_Out, channel2_Kernel42_Valid_Out, channel3_Kernel42_Valid_Out, channel4_Kernel42_Valid_Out, channel5_Kernel42_Valid_Out, channel6_Kernel42_Valid_Out, channel7_Kernel42_Valid_Out, channel8_Kernel42_Valid_Out, channel9_Kernel42_Valid_Out, channel10_Kernel42_Valid_Out, channel11_Kernel42_Valid_Out, channel12_Kernel42_Valid_Out, channel13_Kernel42_Valid_Out, channel14_Kernel42_Valid_Out, channel15_Kernel42_Valid_Out, channel16_Kernel42_Valid_Out, channel17_Kernel42_Valid_Out, channel18_Kernel42_Valid_Out, channel19_Kernel42_Valid_Out, channel20_Kernel42_Valid_Out, channel21_Kernel42_Valid_Out, channel22_Kernel42_Valid_Out, channel23_Kernel42_Valid_Out, channel24_Kernel42_Valid_Out, channel25_Kernel42_Valid_Out, channel26_Kernel42_Valid_Out, channel27_Kernel42_Valid_Out, channel28_Kernel42_Valid_Out, channel29_Kernel42_Valid_Out, channel30_Kernel42_Valid_Out, channel31_Kernel42_Valid_Out, channel32_Kernel42_Valid_Out, channel33_Kernel42_Valid_Out, channel34_Kernel42_Valid_Out, channel35_Kernel42_Valid_Out, channel36_Kernel42_Valid_Out, channel37_Kernel42_Valid_Out, channel38_Kernel42_Valid_Out, channel39_Kernel42_Valid_Out, channel40_Kernel42_Valid_Out, channel41_Kernel42_Valid_Out, channel42_Kernel42_Valid_Out, channel43_Kernel42_Valid_Out, channel44_Kernel42_Valid_Out, channel45_Kernel42_Valid_Out, channel46_Kernel42_Valid_Out, channel47_Kernel42_Valid_Out, channel48_Kernel42_Valid_Out, channel49_Kernel42_Valid_Out, channel50_Kernel42_Valid_Out, channel51_Kernel42_Valid_Out, channel52_Kernel42_Valid_Out, channel53_Kernel42_Valid_Out, channel54_Kernel42_Valid_Out, channel55_Kernel42_Valid_Out, channel56_Kernel42_Valid_Out, channel57_Kernel42_Valid_Out, channel58_Kernel42_Valid_Out, channel59_Kernel42_Valid_Out, channel60_Kernel42_Valid_Out, channel61_Kernel42_Valid_Out, channel62_Kernel42_Valid_Out, channel63_Kernel42_Valid_Out, channel64_Kernel42_Valid_Out;

	assign add_kernel42=channel1_Kernel42_Valid_Out & channel2_Kernel42_Valid_Out & channel3_Kernel42_Valid_Out & channel4_Kernel42_Valid_Out & channel5_Kernel42_Valid_Out & channel6_Kernel42_Valid_Out & channel7_Kernel42_Valid_Out & channel8_Kernel42_Valid_Out & channel9_Kernel42_Valid_Out & channel10_Kernel42_Valid_Out & channel11_Kernel42_Valid_Out & channel12_Kernel42_Valid_Out & channel13_Kernel42_Valid_Out & channel14_Kernel42_Valid_Out & channel15_Kernel42_Valid_Out & channel16_Kernel42_Valid_Out & channel17_Kernel42_Valid_Out & channel18_Kernel42_Valid_Out & channel19_Kernel42_Valid_Out & channel20_Kernel42_Valid_Out & channel21_Kernel42_Valid_Out & channel22_Kernel42_Valid_Out & channel23_Kernel42_Valid_Out & channel24_Kernel42_Valid_Out & channel25_Kernel42_Valid_Out & channel26_Kernel42_Valid_Out & channel27_Kernel42_Valid_Out & channel28_Kernel42_Valid_Out & channel29_Kernel42_Valid_Out & channel30_Kernel42_Valid_Out & channel31_Kernel42_Valid_Out & channel32_Kernel42_Valid_Out & channel33_Kernel42_Valid_Out & channel34_Kernel42_Valid_Out & channel35_Kernel42_Valid_Out & channel36_Kernel42_Valid_Out & channel37_Kernel42_Valid_Out & channel38_Kernel42_Valid_Out & channel39_Kernel42_Valid_Out & channel40_Kernel42_Valid_Out & channel41_Kernel42_Valid_Out & channel42_Kernel42_Valid_Out & channel43_Kernel42_Valid_Out & channel44_Kernel42_Valid_Out & channel45_Kernel42_Valid_Out & channel46_Kernel42_Valid_Out & channel47_Kernel42_Valid_Out & channel48_Kernel42_Valid_Out & channel49_Kernel42_Valid_Out & channel50_Kernel42_Valid_Out & channel51_Kernel42_Valid_Out & channel52_Kernel42_Valid_Out & channel53_Kernel42_Valid_Out & channel54_Kernel42_Valid_Out & channel55_Kernel42_Valid_Out & channel56_Kernel42_Valid_Out & channel57_Kernel42_Valid_Out & channel58_Kernel42_Valid_Out & channel59_Kernel42_Valid_Out & channel60_Kernel42_Valid_Out & channel61_Kernel42_Valid_Out & channel62_Kernel42_Valid_Out & channel63_Kernel42_Valid_Out & channel64_Kernel42_Valid_Out;

	wire channel1_Kernel43_Valid_Out, channel2_Kernel43_Valid_Out, channel3_Kernel43_Valid_Out, channel4_Kernel43_Valid_Out, channel5_Kernel43_Valid_Out, channel6_Kernel43_Valid_Out, channel7_Kernel43_Valid_Out, channel8_Kernel43_Valid_Out, channel9_Kernel43_Valid_Out, channel10_Kernel43_Valid_Out, channel11_Kernel43_Valid_Out, channel12_Kernel43_Valid_Out, channel13_Kernel43_Valid_Out, channel14_Kernel43_Valid_Out, channel15_Kernel43_Valid_Out, channel16_Kernel43_Valid_Out, channel17_Kernel43_Valid_Out, channel18_Kernel43_Valid_Out, channel19_Kernel43_Valid_Out, channel20_Kernel43_Valid_Out, channel21_Kernel43_Valid_Out, channel22_Kernel43_Valid_Out, channel23_Kernel43_Valid_Out, channel24_Kernel43_Valid_Out, channel25_Kernel43_Valid_Out, channel26_Kernel43_Valid_Out, channel27_Kernel43_Valid_Out, channel28_Kernel43_Valid_Out, channel29_Kernel43_Valid_Out, channel30_Kernel43_Valid_Out, channel31_Kernel43_Valid_Out, channel32_Kernel43_Valid_Out, channel33_Kernel43_Valid_Out, channel34_Kernel43_Valid_Out, channel35_Kernel43_Valid_Out, channel36_Kernel43_Valid_Out, channel37_Kernel43_Valid_Out, channel38_Kernel43_Valid_Out, channel39_Kernel43_Valid_Out, channel40_Kernel43_Valid_Out, channel41_Kernel43_Valid_Out, channel42_Kernel43_Valid_Out, channel43_Kernel43_Valid_Out, channel44_Kernel43_Valid_Out, channel45_Kernel43_Valid_Out, channel46_Kernel43_Valid_Out, channel47_Kernel43_Valid_Out, channel48_Kernel43_Valid_Out, channel49_Kernel43_Valid_Out, channel50_Kernel43_Valid_Out, channel51_Kernel43_Valid_Out, channel52_Kernel43_Valid_Out, channel53_Kernel43_Valid_Out, channel54_Kernel43_Valid_Out, channel55_Kernel43_Valid_Out, channel56_Kernel43_Valid_Out, channel57_Kernel43_Valid_Out, channel58_Kernel43_Valid_Out, channel59_Kernel43_Valid_Out, channel60_Kernel43_Valid_Out, channel61_Kernel43_Valid_Out, channel62_Kernel43_Valid_Out, channel63_Kernel43_Valid_Out, channel64_Kernel43_Valid_Out;

	assign add_kernel43=channel1_Kernel43_Valid_Out & channel2_Kernel43_Valid_Out & channel3_Kernel43_Valid_Out & channel4_Kernel43_Valid_Out & channel5_Kernel43_Valid_Out & channel6_Kernel43_Valid_Out & channel7_Kernel43_Valid_Out & channel8_Kernel43_Valid_Out & channel9_Kernel43_Valid_Out & channel10_Kernel43_Valid_Out & channel11_Kernel43_Valid_Out & channel12_Kernel43_Valid_Out & channel13_Kernel43_Valid_Out & channel14_Kernel43_Valid_Out & channel15_Kernel43_Valid_Out & channel16_Kernel43_Valid_Out & channel17_Kernel43_Valid_Out & channel18_Kernel43_Valid_Out & channel19_Kernel43_Valid_Out & channel20_Kernel43_Valid_Out & channel21_Kernel43_Valid_Out & channel22_Kernel43_Valid_Out & channel23_Kernel43_Valid_Out & channel24_Kernel43_Valid_Out & channel25_Kernel43_Valid_Out & channel26_Kernel43_Valid_Out & channel27_Kernel43_Valid_Out & channel28_Kernel43_Valid_Out & channel29_Kernel43_Valid_Out & channel30_Kernel43_Valid_Out & channel31_Kernel43_Valid_Out & channel32_Kernel43_Valid_Out & channel33_Kernel43_Valid_Out & channel34_Kernel43_Valid_Out & channel35_Kernel43_Valid_Out & channel36_Kernel43_Valid_Out & channel37_Kernel43_Valid_Out & channel38_Kernel43_Valid_Out & channel39_Kernel43_Valid_Out & channel40_Kernel43_Valid_Out & channel41_Kernel43_Valid_Out & channel42_Kernel43_Valid_Out & channel43_Kernel43_Valid_Out & channel44_Kernel43_Valid_Out & channel45_Kernel43_Valid_Out & channel46_Kernel43_Valid_Out & channel47_Kernel43_Valid_Out & channel48_Kernel43_Valid_Out & channel49_Kernel43_Valid_Out & channel50_Kernel43_Valid_Out & channel51_Kernel43_Valid_Out & channel52_Kernel43_Valid_Out & channel53_Kernel43_Valid_Out & channel54_Kernel43_Valid_Out & channel55_Kernel43_Valid_Out & channel56_Kernel43_Valid_Out & channel57_Kernel43_Valid_Out & channel58_Kernel43_Valid_Out & channel59_Kernel43_Valid_Out & channel60_Kernel43_Valid_Out & channel61_Kernel43_Valid_Out & channel62_Kernel43_Valid_Out & channel63_Kernel43_Valid_Out & channel64_Kernel43_Valid_Out;

	wire channel1_Kernel44_Valid_Out, channel2_Kernel44_Valid_Out, channel3_Kernel44_Valid_Out, channel4_Kernel44_Valid_Out, channel5_Kernel44_Valid_Out, channel6_Kernel44_Valid_Out, channel7_Kernel44_Valid_Out, channel8_Kernel44_Valid_Out, channel9_Kernel44_Valid_Out, channel10_Kernel44_Valid_Out, channel11_Kernel44_Valid_Out, channel12_Kernel44_Valid_Out, channel13_Kernel44_Valid_Out, channel14_Kernel44_Valid_Out, channel15_Kernel44_Valid_Out, channel16_Kernel44_Valid_Out, channel17_Kernel44_Valid_Out, channel18_Kernel44_Valid_Out, channel19_Kernel44_Valid_Out, channel20_Kernel44_Valid_Out, channel21_Kernel44_Valid_Out, channel22_Kernel44_Valid_Out, channel23_Kernel44_Valid_Out, channel24_Kernel44_Valid_Out, channel25_Kernel44_Valid_Out, channel26_Kernel44_Valid_Out, channel27_Kernel44_Valid_Out, channel28_Kernel44_Valid_Out, channel29_Kernel44_Valid_Out, channel30_Kernel44_Valid_Out, channel31_Kernel44_Valid_Out, channel32_Kernel44_Valid_Out, channel33_Kernel44_Valid_Out, channel34_Kernel44_Valid_Out, channel35_Kernel44_Valid_Out, channel36_Kernel44_Valid_Out, channel37_Kernel44_Valid_Out, channel38_Kernel44_Valid_Out, channel39_Kernel44_Valid_Out, channel40_Kernel44_Valid_Out, channel41_Kernel44_Valid_Out, channel42_Kernel44_Valid_Out, channel43_Kernel44_Valid_Out, channel44_Kernel44_Valid_Out, channel45_Kernel44_Valid_Out, channel46_Kernel44_Valid_Out, channel47_Kernel44_Valid_Out, channel48_Kernel44_Valid_Out, channel49_Kernel44_Valid_Out, channel50_Kernel44_Valid_Out, channel51_Kernel44_Valid_Out, channel52_Kernel44_Valid_Out, channel53_Kernel44_Valid_Out, channel54_Kernel44_Valid_Out, channel55_Kernel44_Valid_Out, channel56_Kernel44_Valid_Out, channel57_Kernel44_Valid_Out, channel58_Kernel44_Valid_Out, channel59_Kernel44_Valid_Out, channel60_Kernel44_Valid_Out, channel61_Kernel44_Valid_Out, channel62_Kernel44_Valid_Out, channel63_Kernel44_Valid_Out, channel64_Kernel44_Valid_Out;

	assign add_kernel44=channel1_Kernel44_Valid_Out & channel2_Kernel44_Valid_Out & channel3_Kernel44_Valid_Out & channel4_Kernel44_Valid_Out & channel5_Kernel44_Valid_Out & channel6_Kernel44_Valid_Out & channel7_Kernel44_Valid_Out & channel8_Kernel44_Valid_Out & channel9_Kernel44_Valid_Out & channel10_Kernel44_Valid_Out & channel11_Kernel44_Valid_Out & channel12_Kernel44_Valid_Out & channel13_Kernel44_Valid_Out & channel14_Kernel44_Valid_Out & channel15_Kernel44_Valid_Out & channel16_Kernel44_Valid_Out & channel17_Kernel44_Valid_Out & channel18_Kernel44_Valid_Out & channel19_Kernel44_Valid_Out & channel20_Kernel44_Valid_Out & channel21_Kernel44_Valid_Out & channel22_Kernel44_Valid_Out & channel23_Kernel44_Valid_Out & channel24_Kernel44_Valid_Out & channel25_Kernel44_Valid_Out & channel26_Kernel44_Valid_Out & channel27_Kernel44_Valid_Out & channel28_Kernel44_Valid_Out & channel29_Kernel44_Valid_Out & channel30_Kernel44_Valid_Out & channel31_Kernel44_Valid_Out & channel32_Kernel44_Valid_Out & channel33_Kernel44_Valid_Out & channel34_Kernel44_Valid_Out & channel35_Kernel44_Valid_Out & channel36_Kernel44_Valid_Out & channel37_Kernel44_Valid_Out & channel38_Kernel44_Valid_Out & channel39_Kernel44_Valid_Out & channel40_Kernel44_Valid_Out & channel41_Kernel44_Valid_Out & channel42_Kernel44_Valid_Out & channel43_Kernel44_Valid_Out & channel44_Kernel44_Valid_Out & channel45_Kernel44_Valid_Out & channel46_Kernel44_Valid_Out & channel47_Kernel44_Valid_Out & channel48_Kernel44_Valid_Out & channel49_Kernel44_Valid_Out & channel50_Kernel44_Valid_Out & channel51_Kernel44_Valid_Out & channel52_Kernel44_Valid_Out & channel53_Kernel44_Valid_Out & channel54_Kernel44_Valid_Out & channel55_Kernel44_Valid_Out & channel56_Kernel44_Valid_Out & channel57_Kernel44_Valid_Out & channel58_Kernel44_Valid_Out & channel59_Kernel44_Valid_Out & channel60_Kernel44_Valid_Out & channel61_Kernel44_Valid_Out & channel62_Kernel44_Valid_Out & channel63_Kernel44_Valid_Out & channel64_Kernel44_Valid_Out;

	wire channel1_Kernel45_Valid_Out, channel2_Kernel45_Valid_Out, channel3_Kernel45_Valid_Out, channel4_Kernel45_Valid_Out, channel5_Kernel45_Valid_Out, channel6_Kernel45_Valid_Out, channel7_Kernel45_Valid_Out, channel8_Kernel45_Valid_Out, channel9_Kernel45_Valid_Out, channel10_Kernel45_Valid_Out, channel11_Kernel45_Valid_Out, channel12_Kernel45_Valid_Out, channel13_Kernel45_Valid_Out, channel14_Kernel45_Valid_Out, channel15_Kernel45_Valid_Out, channel16_Kernel45_Valid_Out, channel17_Kernel45_Valid_Out, channel18_Kernel45_Valid_Out, channel19_Kernel45_Valid_Out, channel20_Kernel45_Valid_Out, channel21_Kernel45_Valid_Out, channel22_Kernel45_Valid_Out, channel23_Kernel45_Valid_Out, channel24_Kernel45_Valid_Out, channel25_Kernel45_Valid_Out, channel26_Kernel45_Valid_Out, channel27_Kernel45_Valid_Out, channel28_Kernel45_Valid_Out, channel29_Kernel45_Valid_Out, channel30_Kernel45_Valid_Out, channel31_Kernel45_Valid_Out, channel32_Kernel45_Valid_Out, channel33_Kernel45_Valid_Out, channel34_Kernel45_Valid_Out, channel35_Kernel45_Valid_Out, channel36_Kernel45_Valid_Out, channel37_Kernel45_Valid_Out, channel38_Kernel45_Valid_Out, channel39_Kernel45_Valid_Out, channel40_Kernel45_Valid_Out, channel41_Kernel45_Valid_Out, channel42_Kernel45_Valid_Out, channel43_Kernel45_Valid_Out, channel44_Kernel45_Valid_Out, channel45_Kernel45_Valid_Out, channel46_Kernel45_Valid_Out, channel47_Kernel45_Valid_Out, channel48_Kernel45_Valid_Out, channel49_Kernel45_Valid_Out, channel50_Kernel45_Valid_Out, channel51_Kernel45_Valid_Out, channel52_Kernel45_Valid_Out, channel53_Kernel45_Valid_Out, channel54_Kernel45_Valid_Out, channel55_Kernel45_Valid_Out, channel56_Kernel45_Valid_Out, channel57_Kernel45_Valid_Out, channel58_Kernel45_Valid_Out, channel59_Kernel45_Valid_Out, channel60_Kernel45_Valid_Out, channel61_Kernel45_Valid_Out, channel62_Kernel45_Valid_Out, channel63_Kernel45_Valid_Out, channel64_Kernel45_Valid_Out;

	assign add_kernel45=channel1_Kernel45_Valid_Out & channel2_Kernel45_Valid_Out & channel3_Kernel45_Valid_Out & channel4_Kernel45_Valid_Out & channel5_Kernel45_Valid_Out & channel6_Kernel45_Valid_Out & channel7_Kernel45_Valid_Out & channel8_Kernel45_Valid_Out & channel9_Kernel45_Valid_Out & channel10_Kernel45_Valid_Out & channel11_Kernel45_Valid_Out & channel12_Kernel45_Valid_Out & channel13_Kernel45_Valid_Out & channel14_Kernel45_Valid_Out & channel15_Kernel45_Valid_Out & channel16_Kernel45_Valid_Out & channel17_Kernel45_Valid_Out & channel18_Kernel45_Valid_Out & channel19_Kernel45_Valid_Out & channel20_Kernel45_Valid_Out & channel21_Kernel45_Valid_Out & channel22_Kernel45_Valid_Out & channel23_Kernel45_Valid_Out & channel24_Kernel45_Valid_Out & channel25_Kernel45_Valid_Out & channel26_Kernel45_Valid_Out & channel27_Kernel45_Valid_Out & channel28_Kernel45_Valid_Out & channel29_Kernel45_Valid_Out & channel30_Kernel45_Valid_Out & channel31_Kernel45_Valid_Out & channel32_Kernel45_Valid_Out & channel33_Kernel45_Valid_Out & channel34_Kernel45_Valid_Out & channel35_Kernel45_Valid_Out & channel36_Kernel45_Valid_Out & channel37_Kernel45_Valid_Out & channel38_Kernel45_Valid_Out & channel39_Kernel45_Valid_Out & channel40_Kernel45_Valid_Out & channel41_Kernel45_Valid_Out & channel42_Kernel45_Valid_Out & channel43_Kernel45_Valid_Out & channel44_Kernel45_Valid_Out & channel45_Kernel45_Valid_Out & channel46_Kernel45_Valid_Out & channel47_Kernel45_Valid_Out & channel48_Kernel45_Valid_Out & channel49_Kernel45_Valid_Out & channel50_Kernel45_Valid_Out & channel51_Kernel45_Valid_Out & channel52_Kernel45_Valid_Out & channel53_Kernel45_Valid_Out & channel54_Kernel45_Valid_Out & channel55_Kernel45_Valid_Out & channel56_Kernel45_Valid_Out & channel57_Kernel45_Valid_Out & channel58_Kernel45_Valid_Out & channel59_Kernel45_Valid_Out & channel60_Kernel45_Valid_Out & channel61_Kernel45_Valid_Out & channel62_Kernel45_Valid_Out & channel63_Kernel45_Valid_Out & channel64_Kernel45_Valid_Out;

	wire channel1_Kernel46_Valid_Out, channel2_Kernel46_Valid_Out, channel3_Kernel46_Valid_Out, channel4_Kernel46_Valid_Out, channel5_Kernel46_Valid_Out, channel6_Kernel46_Valid_Out, channel7_Kernel46_Valid_Out, channel8_Kernel46_Valid_Out, channel9_Kernel46_Valid_Out, channel10_Kernel46_Valid_Out, channel11_Kernel46_Valid_Out, channel12_Kernel46_Valid_Out, channel13_Kernel46_Valid_Out, channel14_Kernel46_Valid_Out, channel15_Kernel46_Valid_Out, channel16_Kernel46_Valid_Out, channel17_Kernel46_Valid_Out, channel18_Kernel46_Valid_Out, channel19_Kernel46_Valid_Out, channel20_Kernel46_Valid_Out, channel21_Kernel46_Valid_Out, channel22_Kernel46_Valid_Out, channel23_Kernel46_Valid_Out, channel24_Kernel46_Valid_Out, channel25_Kernel46_Valid_Out, channel26_Kernel46_Valid_Out, channel27_Kernel46_Valid_Out, channel28_Kernel46_Valid_Out, channel29_Kernel46_Valid_Out, channel30_Kernel46_Valid_Out, channel31_Kernel46_Valid_Out, channel32_Kernel46_Valid_Out, channel33_Kernel46_Valid_Out, channel34_Kernel46_Valid_Out, channel35_Kernel46_Valid_Out, channel36_Kernel46_Valid_Out, channel37_Kernel46_Valid_Out, channel38_Kernel46_Valid_Out, channel39_Kernel46_Valid_Out, channel40_Kernel46_Valid_Out, channel41_Kernel46_Valid_Out, channel42_Kernel46_Valid_Out, channel43_Kernel46_Valid_Out, channel44_Kernel46_Valid_Out, channel45_Kernel46_Valid_Out, channel46_Kernel46_Valid_Out, channel47_Kernel46_Valid_Out, channel48_Kernel46_Valid_Out, channel49_Kernel46_Valid_Out, channel50_Kernel46_Valid_Out, channel51_Kernel46_Valid_Out, channel52_Kernel46_Valid_Out, channel53_Kernel46_Valid_Out, channel54_Kernel46_Valid_Out, channel55_Kernel46_Valid_Out, channel56_Kernel46_Valid_Out, channel57_Kernel46_Valid_Out, channel58_Kernel46_Valid_Out, channel59_Kernel46_Valid_Out, channel60_Kernel46_Valid_Out, channel61_Kernel46_Valid_Out, channel62_Kernel46_Valid_Out, channel63_Kernel46_Valid_Out, channel64_Kernel46_Valid_Out;

	assign add_kernel46=channel1_Kernel46_Valid_Out & channel2_Kernel46_Valid_Out & channel3_Kernel46_Valid_Out & channel4_Kernel46_Valid_Out & channel5_Kernel46_Valid_Out & channel6_Kernel46_Valid_Out & channel7_Kernel46_Valid_Out & channel8_Kernel46_Valid_Out & channel9_Kernel46_Valid_Out & channel10_Kernel46_Valid_Out & channel11_Kernel46_Valid_Out & channel12_Kernel46_Valid_Out & channel13_Kernel46_Valid_Out & channel14_Kernel46_Valid_Out & channel15_Kernel46_Valid_Out & channel16_Kernel46_Valid_Out & channel17_Kernel46_Valid_Out & channel18_Kernel46_Valid_Out & channel19_Kernel46_Valid_Out & channel20_Kernel46_Valid_Out & channel21_Kernel46_Valid_Out & channel22_Kernel46_Valid_Out & channel23_Kernel46_Valid_Out & channel24_Kernel46_Valid_Out & channel25_Kernel46_Valid_Out & channel26_Kernel46_Valid_Out & channel27_Kernel46_Valid_Out & channel28_Kernel46_Valid_Out & channel29_Kernel46_Valid_Out & channel30_Kernel46_Valid_Out & channel31_Kernel46_Valid_Out & channel32_Kernel46_Valid_Out & channel33_Kernel46_Valid_Out & channel34_Kernel46_Valid_Out & channel35_Kernel46_Valid_Out & channel36_Kernel46_Valid_Out & channel37_Kernel46_Valid_Out & channel38_Kernel46_Valid_Out & channel39_Kernel46_Valid_Out & channel40_Kernel46_Valid_Out & channel41_Kernel46_Valid_Out & channel42_Kernel46_Valid_Out & channel43_Kernel46_Valid_Out & channel44_Kernel46_Valid_Out & channel45_Kernel46_Valid_Out & channel46_Kernel46_Valid_Out & channel47_Kernel46_Valid_Out & channel48_Kernel46_Valid_Out & channel49_Kernel46_Valid_Out & channel50_Kernel46_Valid_Out & channel51_Kernel46_Valid_Out & channel52_Kernel46_Valid_Out & channel53_Kernel46_Valid_Out & channel54_Kernel46_Valid_Out & channel55_Kernel46_Valid_Out & channel56_Kernel46_Valid_Out & channel57_Kernel46_Valid_Out & channel58_Kernel46_Valid_Out & channel59_Kernel46_Valid_Out & channel60_Kernel46_Valid_Out & channel61_Kernel46_Valid_Out & channel62_Kernel46_Valid_Out & channel63_Kernel46_Valid_Out & channel64_Kernel46_Valid_Out;

	wire channel1_Kernel47_Valid_Out, channel2_Kernel47_Valid_Out, channel3_Kernel47_Valid_Out, channel4_Kernel47_Valid_Out, channel5_Kernel47_Valid_Out, channel6_Kernel47_Valid_Out, channel7_Kernel47_Valid_Out, channel8_Kernel47_Valid_Out, channel9_Kernel47_Valid_Out, channel10_Kernel47_Valid_Out, channel11_Kernel47_Valid_Out, channel12_Kernel47_Valid_Out, channel13_Kernel47_Valid_Out, channel14_Kernel47_Valid_Out, channel15_Kernel47_Valid_Out, channel16_Kernel47_Valid_Out, channel17_Kernel47_Valid_Out, channel18_Kernel47_Valid_Out, channel19_Kernel47_Valid_Out, channel20_Kernel47_Valid_Out, channel21_Kernel47_Valid_Out, channel22_Kernel47_Valid_Out, channel23_Kernel47_Valid_Out, channel24_Kernel47_Valid_Out, channel25_Kernel47_Valid_Out, channel26_Kernel47_Valid_Out, channel27_Kernel47_Valid_Out, channel28_Kernel47_Valid_Out, channel29_Kernel47_Valid_Out, channel30_Kernel47_Valid_Out, channel31_Kernel47_Valid_Out, channel32_Kernel47_Valid_Out, channel33_Kernel47_Valid_Out, channel34_Kernel47_Valid_Out, channel35_Kernel47_Valid_Out, channel36_Kernel47_Valid_Out, channel37_Kernel47_Valid_Out, channel38_Kernel47_Valid_Out, channel39_Kernel47_Valid_Out, channel40_Kernel47_Valid_Out, channel41_Kernel47_Valid_Out, channel42_Kernel47_Valid_Out, channel43_Kernel47_Valid_Out, channel44_Kernel47_Valid_Out, channel45_Kernel47_Valid_Out, channel46_Kernel47_Valid_Out, channel47_Kernel47_Valid_Out, channel48_Kernel47_Valid_Out, channel49_Kernel47_Valid_Out, channel50_Kernel47_Valid_Out, channel51_Kernel47_Valid_Out, channel52_Kernel47_Valid_Out, channel53_Kernel47_Valid_Out, channel54_Kernel47_Valid_Out, channel55_Kernel47_Valid_Out, channel56_Kernel47_Valid_Out, channel57_Kernel47_Valid_Out, channel58_Kernel47_Valid_Out, channel59_Kernel47_Valid_Out, channel60_Kernel47_Valid_Out, channel61_Kernel47_Valid_Out, channel62_Kernel47_Valid_Out, channel63_Kernel47_Valid_Out, channel64_Kernel47_Valid_Out;

	assign add_kernel47=channel1_Kernel47_Valid_Out & channel2_Kernel47_Valid_Out & channel3_Kernel47_Valid_Out & channel4_Kernel47_Valid_Out & channel5_Kernel47_Valid_Out & channel6_Kernel47_Valid_Out & channel7_Kernel47_Valid_Out & channel8_Kernel47_Valid_Out & channel9_Kernel47_Valid_Out & channel10_Kernel47_Valid_Out & channel11_Kernel47_Valid_Out & channel12_Kernel47_Valid_Out & channel13_Kernel47_Valid_Out & channel14_Kernel47_Valid_Out & channel15_Kernel47_Valid_Out & channel16_Kernel47_Valid_Out & channel17_Kernel47_Valid_Out & channel18_Kernel47_Valid_Out & channel19_Kernel47_Valid_Out & channel20_Kernel47_Valid_Out & channel21_Kernel47_Valid_Out & channel22_Kernel47_Valid_Out & channel23_Kernel47_Valid_Out & channel24_Kernel47_Valid_Out & channel25_Kernel47_Valid_Out & channel26_Kernel47_Valid_Out & channel27_Kernel47_Valid_Out & channel28_Kernel47_Valid_Out & channel29_Kernel47_Valid_Out & channel30_Kernel47_Valid_Out & channel31_Kernel47_Valid_Out & channel32_Kernel47_Valid_Out & channel33_Kernel47_Valid_Out & channel34_Kernel47_Valid_Out & channel35_Kernel47_Valid_Out & channel36_Kernel47_Valid_Out & channel37_Kernel47_Valid_Out & channel38_Kernel47_Valid_Out & channel39_Kernel47_Valid_Out & channel40_Kernel47_Valid_Out & channel41_Kernel47_Valid_Out & channel42_Kernel47_Valid_Out & channel43_Kernel47_Valid_Out & channel44_Kernel47_Valid_Out & channel45_Kernel47_Valid_Out & channel46_Kernel47_Valid_Out & channel47_Kernel47_Valid_Out & channel48_Kernel47_Valid_Out & channel49_Kernel47_Valid_Out & channel50_Kernel47_Valid_Out & channel51_Kernel47_Valid_Out & channel52_Kernel47_Valid_Out & channel53_Kernel47_Valid_Out & channel54_Kernel47_Valid_Out & channel55_Kernel47_Valid_Out & channel56_Kernel47_Valid_Out & channel57_Kernel47_Valid_Out & channel58_Kernel47_Valid_Out & channel59_Kernel47_Valid_Out & channel60_Kernel47_Valid_Out & channel61_Kernel47_Valid_Out & channel62_Kernel47_Valid_Out & channel63_Kernel47_Valid_Out & channel64_Kernel47_Valid_Out;

	wire channel1_Kernel48_Valid_Out, channel2_Kernel48_Valid_Out, channel3_Kernel48_Valid_Out, channel4_Kernel48_Valid_Out, channel5_Kernel48_Valid_Out, channel6_Kernel48_Valid_Out, channel7_Kernel48_Valid_Out, channel8_Kernel48_Valid_Out, channel9_Kernel48_Valid_Out, channel10_Kernel48_Valid_Out, channel11_Kernel48_Valid_Out, channel12_Kernel48_Valid_Out, channel13_Kernel48_Valid_Out, channel14_Kernel48_Valid_Out, channel15_Kernel48_Valid_Out, channel16_Kernel48_Valid_Out, channel17_Kernel48_Valid_Out, channel18_Kernel48_Valid_Out, channel19_Kernel48_Valid_Out, channel20_Kernel48_Valid_Out, channel21_Kernel48_Valid_Out, channel22_Kernel48_Valid_Out, channel23_Kernel48_Valid_Out, channel24_Kernel48_Valid_Out, channel25_Kernel48_Valid_Out, channel26_Kernel48_Valid_Out, channel27_Kernel48_Valid_Out, channel28_Kernel48_Valid_Out, channel29_Kernel48_Valid_Out, channel30_Kernel48_Valid_Out, channel31_Kernel48_Valid_Out, channel32_Kernel48_Valid_Out, channel33_Kernel48_Valid_Out, channel34_Kernel48_Valid_Out, channel35_Kernel48_Valid_Out, channel36_Kernel48_Valid_Out, channel37_Kernel48_Valid_Out, channel38_Kernel48_Valid_Out, channel39_Kernel48_Valid_Out, channel40_Kernel48_Valid_Out, channel41_Kernel48_Valid_Out, channel42_Kernel48_Valid_Out, channel43_Kernel48_Valid_Out, channel44_Kernel48_Valid_Out, channel45_Kernel48_Valid_Out, channel46_Kernel48_Valid_Out, channel47_Kernel48_Valid_Out, channel48_Kernel48_Valid_Out, channel49_Kernel48_Valid_Out, channel50_Kernel48_Valid_Out, channel51_Kernel48_Valid_Out, channel52_Kernel48_Valid_Out, channel53_Kernel48_Valid_Out, channel54_Kernel48_Valid_Out, channel55_Kernel48_Valid_Out, channel56_Kernel48_Valid_Out, channel57_Kernel48_Valid_Out, channel58_Kernel48_Valid_Out, channel59_Kernel48_Valid_Out, channel60_Kernel48_Valid_Out, channel61_Kernel48_Valid_Out, channel62_Kernel48_Valid_Out, channel63_Kernel48_Valid_Out, channel64_Kernel48_Valid_Out;

	assign add_kernel48=channel1_Kernel48_Valid_Out & channel2_Kernel48_Valid_Out & channel3_Kernel48_Valid_Out & channel4_Kernel48_Valid_Out & channel5_Kernel48_Valid_Out & channel6_Kernel48_Valid_Out & channel7_Kernel48_Valid_Out & channel8_Kernel48_Valid_Out & channel9_Kernel48_Valid_Out & channel10_Kernel48_Valid_Out & channel11_Kernel48_Valid_Out & channel12_Kernel48_Valid_Out & channel13_Kernel48_Valid_Out & channel14_Kernel48_Valid_Out & channel15_Kernel48_Valid_Out & channel16_Kernel48_Valid_Out & channel17_Kernel48_Valid_Out & channel18_Kernel48_Valid_Out & channel19_Kernel48_Valid_Out & channel20_Kernel48_Valid_Out & channel21_Kernel48_Valid_Out & channel22_Kernel48_Valid_Out & channel23_Kernel48_Valid_Out & channel24_Kernel48_Valid_Out & channel25_Kernel48_Valid_Out & channel26_Kernel48_Valid_Out & channel27_Kernel48_Valid_Out & channel28_Kernel48_Valid_Out & channel29_Kernel48_Valid_Out & channel30_Kernel48_Valid_Out & channel31_Kernel48_Valid_Out & channel32_Kernel48_Valid_Out & channel33_Kernel48_Valid_Out & channel34_Kernel48_Valid_Out & channel35_Kernel48_Valid_Out & channel36_Kernel48_Valid_Out & channel37_Kernel48_Valid_Out & channel38_Kernel48_Valid_Out & channel39_Kernel48_Valid_Out & channel40_Kernel48_Valid_Out & channel41_Kernel48_Valid_Out & channel42_Kernel48_Valid_Out & channel43_Kernel48_Valid_Out & channel44_Kernel48_Valid_Out & channel45_Kernel48_Valid_Out & channel46_Kernel48_Valid_Out & channel47_Kernel48_Valid_Out & channel48_Kernel48_Valid_Out & channel49_Kernel48_Valid_Out & channel50_Kernel48_Valid_Out & channel51_Kernel48_Valid_Out & channel52_Kernel48_Valid_Out & channel53_Kernel48_Valid_Out & channel54_Kernel48_Valid_Out & channel55_Kernel48_Valid_Out & channel56_Kernel48_Valid_Out & channel57_Kernel48_Valid_Out & channel58_Kernel48_Valid_Out & channel59_Kernel48_Valid_Out & channel60_Kernel48_Valid_Out & channel61_Kernel48_Valid_Out & channel62_Kernel48_Valid_Out & channel63_Kernel48_Valid_Out & channel64_Kernel48_Valid_Out;

	wire channel1_Kernel49_Valid_Out, channel2_Kernel49_Valid_Out, channel3_Kernel49_Valid_Out, channel4_Kernel49_Valid_Out, channel5_Kernel49_Valid_Out, channel6_Kernel49_Valid_Out, channel7_Kernel49_Valid_Out, channel8_Kernel49_Valid_Out, channel9_Kernel49_Valid_Out, channel10_Kernel49_Valid_Out, channel11_Kernel49_Valid_Out, channel12_Kernel49_Valid_Out, channel13_Kernel49_Valid_Out, channel14_Kernel49_Valid_Out, channel15_Kernel49_Valid_Out, channel16_Kernel49_Valid_Out, channel17_Kernel49_Valid_Out, channel18_Kernel49_Valid_Out, channel19_Kernel49_Valid_Out, channel20_Kernel49_Valid_Out, channel21_Kernel49_Valid_Out, channel22_Kernel49_Valid_Out, channel23_Kernel49_Valid_Out, channel24_Kernel49_Valid_Out, channel25_Kernel49_Valid_Out, channel26_Kernel49_Valid_Out, channel27_Kernel49_Valid_Out, channel28_Kernel49_Valid_Out, channel29_Kernel49_Valid_Out, channel30_Kernel49_Valid_Out, channel31_Kernel49_Valid_Out, channel32_Kernel49_Valid_Out, channel33_Kernel49_Valid_Out, channel34_Kernel49_Valid_Out, channel35_Kernel49_Valid_Out, channel36_Kernel49_Valid_Out, channel37_Kernel49_Valid_Out, channel38_Kernel49_Valid_Out, channel39_Kernel49_Valid_Out, channel40_Kernel49_Valid_Out, channel41_Kernel49_Valid_Out, channel42_Kernel49_Valid_Out, channel43_Kernel49_Valid_Out, channel44_Kernel49_Valid_Out, channel45_Kernel49_Valid_Out, channel46_Kernel49_Valid_Out, channel47_Kernel49_Valid_Out, channel48_Kernel49_Valid_Out, channel49_Kernel49_Valid_Out, channel50_Kernel49_Valid_Out, channel51_Kernel49_Valid_Out, channel52_Kernel49_Valid_Out, channel53_Kernel49_Valid_Out, channel54_Kernel49_Valid_Out, channel55_Kernel49_Valid_Out, channel56_Kernel49_Valid_Out, channel57_Kernel49_Valid_Out, channel58_Kernel49_Valid_Out, channel59_Kernel49_Valid_Out, channel60_Kernel49_Valid_Out, channel61_Kernel49_Valid_Out, channel62_Kernel49_Valid_Out, channel63_Kernel49_Valid_Out, channel64_Kernel49_Valid_Out;

	assign add_kernel49=channel1_Kernel49_Valid_Out & channel2_Kernel49_Valid_Out & channel3_Kernel49_Valid_Out & channel4_Kernel49_Valid_Out & channel5_Kernel49_Valid_Out & channel6_Kernel49_Valid_Out & channel7_Kernel49_Valid_Out & channel8_Kernel49_Valid_Out & channel9_Kernel49_Valid_Out & channel10_Kernel49_Valid_Out & channel11_Kernel49_Valid_Out & channel12_Kernel49_Valid_Out & channel13_Kernel49_Valid_Out & channel14_Kernel49_Valid_Out & channel15_Kernel49_Valid_Out & channel16_Kernel49_Valid_Out & channel17_Kernel49_Valid_Out & channel18_Kernel49_Valid_Out & channel19_Kernel49_Valid_Out & channel20_Kernel49_Valid_Out & channel21_Kernel49_Valid_Out & channel22_Kernel49_Valid_Out & channel23_Kernel49_Valid_Out & channel24_Kernel49_Valid_Out & channel25_Kernel49_Valid_Out & channel26_Kernel49_Valid_Out & channel27_Kernel49_Valid_Out & channel28_Kernel49_Valid_Out & channel29_Kernel49_Valid_Out & channel30_Kernel49_Valid_Out & channel31_Kernel49_Valid_Out & channel32_Kernel49_Valid_Out & channel33_Kernel49_Valid_Out & channel34_Kernel49_Valid_Out & channel35_Kernel49_Valid_Out & channel36_Kernel49_Valid_Out & channel37_Kernel49_Valid_Out & channel38_Kernel49_Valid_Out & channel39_Kernel49_Valid_Out & channel40_Kernel49_Valid_Out & channel41_Kernel49_Valid_Out & channel42_Kernel49_Valid_Out & channel43_Kernel49_Valid_Out & channel44_Kernel49_Valid_Out & channel45_Kernel49_Valid_Out & channel46_Kernel49_Valid_Out & channel47_Kernel49_Valid_Out & channel48_Kernel49_Valid_Out & channel49_Kernel49_Valid_Out & channel50_Kernel49_Valid_Out & channel51_Kernel49_Valid_Out & channel52_Kernel49_Valid_Out & channel53_Kernel49_Valid_Out & channel54_Kernel49_Valid_Out & channel55_Kernel49_Valid_Out & channel56_Kernel49_Valid_Out & channel57_Kernel49_Valid_Out & channel58_Kernel49_Valid_Out & channel59_Kernel49_Valid_Out & channel60_Kernel49_Valid_Out & channel61_Kernel49_Valid_Out & channel62_Kernel49_Valid_Out & channel63_Kernel49_Valid_Out & channel64_Kernel49_Valid_Out;

	wire channel1_Kernel50_Valid_Out, channel2_Kernel50_Valid_Out, channel3_Kernel50_Valid_Out, channel4_Kernel50_Valid_Out, channel5_Kernel50_Valid_Out, channel6_Kernel50_Valid_Out, channel7_Kernel50_Valid_Out, channel8_Kernel50_Valid_Out, channel9_Kernel50_Valid_Out, channel10_Kernel50_Valid_Out, channel11_Kernel50_Valid_Out, channel12_Kernel50_Valid_Out, channel13_Kernel50_Valid_Out, channel14_Kernel50_Valid_Out, channel15_Kernel50_Valid_Out, channel16_Kernel50_Valid_Out, channel17_Kernel50_Valid_Out, channel18_Kernel50_Valid_Out, channel19_Kernel50_Valid_Out, channel20_Kernel50_Valid_Out, channel21_Kernel50_Valid_Out, channel22_Kernel50_Valid_Out, channel23_Kernel50_Valid_Out, channel24_Kernel50_Valid_Out, channel25_Kernel50_Valid_Out, channel26_Kernel50_Valid_Out, channel27_Kernel50_Valid_Out, channel28_Kernel50_Valid_Out, channel29_Kernel50_Valid_Out, channel30_Kernel50_Valid_Out, channel31_Kernel50_Valid_Out, channel32_Kernel50_Valid_Out, channel33_Kernel50_Valid_Out, channel34_Kernel50_Valid_Out, channel35_Kernel50_Valid_Out, channel36_Kernel50_Valid_Out, channel37_Kernel50_Valid_Out, channel38_Kernel50_Valid_Out, channel39_Kernel50_Valid_Out, channel40_Kernel50_Valid_Out, channel41_Kernel50_Valid_Out, channel42_Kernel50_Valid_Out, channel43_Kernel50_Valid_Out, channel44_Kernel50_Valid_Out, channel45_Kernel50_Valid_Out, channel46_Kernel50_Valid_Out, channel47_Kernel50_Valid_Out, channel48_Kernel50_Valid_Out, channel49_Kernel50_Valid_Out, channel50_Kernel50_Valid_Out, channel51_Kernel50_Valid_Out, channel52_Kernel50_Valid_Out, channel53_Kernel50_Valid_Out, channel54_Kernel50_Valid_Out, channel55_Kernel50_Valid_Out, channel56_Kernel50_Valid_Out, channel57_Kernel50_Valid_Out, channel58_Kernel50_Valid_Out, channel59_Kernel50_Valid_Out, channel60_Kernel50_Valid_Out, channel61_Kernel50_Valid_Out, channel62_Kernel50_Valid_Out, channel63_Kernel50_Valid_Out, channel64_Kernel50_Valid_Out;

	assign add_kernel50=channel1_Kernel50_Valid_Out & channel2_Kernel50_Valid_Out & channel3_Kernel50_Valid_Out & channel4_Kernel50_Valid_Out & channel5_Kernel50_Valid_Out & channel6_Kernel50_Valid_Out & channel7_Kernel50_Valid_Out & channel8_Kernel50_Valid_Out & channel9_Kernel50_Valid_Out & channel10_Kernel50_Valid_Out & channel11_Kernel50_Valid_Out & channel12_Kernel50_Valid_Out & channel13_Kernel50_Valid_Out & channel14_Kernel50_Valid_Out & channel15_Kernel50_Valid_Out & channel16_Kernel50_Valid_Out & channel17_Kernel50_Valid_Out & channel18_Kernel50_Valid_Out & channel19_Kernel50_Valid_Out & channel20_Kernel50_Valid_Out & channel21_Kernel50_Valid_Out & channel22_Kernel50_Valid_Out & channel23_Kernel50_Valid_Out & channel24_Kernel50_Valid_Out & channel25_Kernel50_Valid_Out & channel26_Kernel50_Valid_Out & channel27_Kernel50_Valid_Out & channel28_Kernel50_Valid_Out & channel29_Kernel50_Valid_Out & channel30_Kernel50_Valid_Out & channel31_Kernel50_Valid_Out & channel32_Kernel50_Valid_Out & channel33_Kernel50_Valid_Out & channel34_Kernel50_Valid_Out & channel35_Kernel50_Valid_Out & channel36_Kernel50_Valid_Out & channel37_Kernel50_Valid_Out & channel38_Kernel50_Valid_Out & channel39_Kernel50_Valid_Out & channel40_Kernel50_Valid_Out & channel41_Kernel50_Valid_Out & channel42_Kernel50_Valid_Out & channel43_Kernel50_Valid_Out & channel44_Kernel50_Valid_Out & channel45_Kernel50_Valid_Out & channel46_Kernel50_Valid_Out & channel47_Kernel50_Valid_Out & channel48_Kernel50_Valid_Out & channel49_Kernel50_Valid_Out & channel50_Kernel50_Valid_Out & channel51_Kernel50_Valid_Out & channel52_Kernel50_Valid_Out & channel53_Kernel50_Valid_Out & channel54_Kernel50_Valid_Out & channel55_Kernel50_Valid_Out & channel56_Kernel50_Valid_Out & channel57_Kernel50_Valid_Out & channel58_Kernel50_Valid_Out & channel59_Kernel50_Valid_Out & channel60_Kernel50_Valid_Out & channel61_Kernel50_Valid_Out & channel62_Kernel50_Valid_Out & channel63_Kernel50_Valid_Out & channel64_Kernel50_Valid_Out;

	wire channel1_Kernel51_Valid_Out, channel2_Kernel51_Valid_Out, channel3_Kernel51_Valid_Out, channel4_Kernel51_Valid_Out, channel5_Kernel51_Valid_Out, channel6_Kernel51_Valid_Out, channel7_Kernel51_Valid_Out, channel8_Kernel51_Valid_Out, channel9_Kernel51_Valid_Out, channel10_Kernel51_Valid_Out, channel11_Kernel51_Valid_Out, channel12_Kernel51_Valid_Out, channel13_Kernel51_Valid_Out, channel14_Kernel51_Valid_Out, channel15_Kernel51_Valid_Out, channel16_Kernel51_Valid_Out, channel17_Kernel51_Valid_Out, channel18_Kernel51_Valid_Out, channel19_Kernel51_Valid_Out, channel20_Kernel51_Valid_Out, channel21_Kernel51_Valid_Out, channel22_Kernel51_Valid_Out, channel23_Kernel51_Valid_Out, channel24_Kernel51_Valid_Out, channel25_Kernel51_Valid_Out, channel26_Kernel51_Valid_Out, channel27_Kernel51_Valid_Out, channel28_Kernel51_Valid_Out, channel29_Kernel51_Valid_Out, channel30_Kernel51_Valid_Out, channel31_Kernel51_Valid_Out, channel32_Kernel51_Valid_Out, channel33_Kernel51_Valid_Out, channel34_Kernel51_Valid_Out, channel35_Kernel51_Valid_Out, channel36_Kernel51_Valid_Out, channel37_Kernel51_Valid_Out, channel38_Kernel51_Valid_Out, channel39_Kernel51_Valid_Out, channel40_Kernel51_Valid_Out, channel41_Kernel51_Valid_Out, channel42_Kernel51_Valid_Out, channel43_Kernel51_Valid_Out, channel44_Kernel51_Valid_Out, channel45_Kernel51_Valid_Out, channel46_Kernel51_Valid_Out, channel47_Kernel51_Valid_Out, channel48_Kernel51_Valid_Out, channel49_Kernel51_Valid_Out, channel50_Kernel51_Valid_Out, channel51_Kernel51_Valid_Out, channel52_Kernel51_Valid_Out, channel53_Kernel51_Valid_Out, channel54_Kernel51_Valid_Out, channel55_Kernel51_Valid_Out, channel56_Kernel51_Valid_Out, channel57_Kernel51_Valid_Out, channel58_Kernel51_Valid_Out, channel59_Kernel51_Valid_Out, channel60_Kernel51_Valid_Out, channel61_Kernel51_Valid_Out, channel62_Kernel51_Valid_Out, channel63_Kernel51_Valid_Out, channel64_Kernel51_Valid_Out;

	assign add_kernel51=channel1_Kernel51_Valid_Out & channel2_Kernel51_Valid_Out & channel3_Kernel51_Valid_Out & channel4_Kernel51_Valid_Out & channel5_Kernel51_Valid_Out & channel6_Kernel51_Valid_Out & channel7_Kernel51_Valid_Out & channel8_Kernel51_Valid_Out & channel9_Kernel51_Valid_Out & channel10_Kernel51_Valid_Out & channel11_Kernel51_Valid_Out & channel12_Kernel51_Valid_Out & channel13_Kernel51_Valid_Out & channel14_Kernel51_Valid_Out & channel15_Kernel51_Valid_Out & channel16_Kernel51_Valid_Out & channel17_Kernel51_Valid_Out & channel18_Kernel51_Valid_Out & channel19_Kernel51_Valid_Out & channel20_Kernel51_Valid_Out & channel21_Kernel51_Valid_Out & channel22_Kernel51_Valid_Out & channel23_Kernel51_Valid_Out & channel24_Kernel51_Valid_Out & channel25_Kernel51_Valid_Out & channel26_Kernel51_Valid_Out & channel27_Kernel51_Valid_Out & channel28_Kernel51_Valid_Out & channel29_Kernel51_Valid_Out & channel30_Kernel51_Valid_Out & channel31_Kernel51_Valid_Out & channel32_Kernel51_Valid_Out & channel33_Kernel51_Valid_Out & channel34_Kernel51_Valid_Out & channel35_Kernel51_Valid_Out & channel36_Kernel51_Valid_Out & channel37_Kernel51_Valid_Out & channel38_Kernel51_Valid_Out & channel39_Kernel51_Valid_Out & channel40_Kernel51_Valid_Out & channel41_Kernel51_Valid_Out & channel42_Kernel51_Valid_Out & channel43_Kernel51_Valid_Out & channel44_Kernel51_Valid_Out & channel45_Kernel51_Valid_Out & channel46_Kernel51_Valid_Out & channel47_Kernel51_Valid_Out & channel48_Kernel51_Valid_Out & channel49_Kernel51_Valid_Out & channel50_Kernel51_Valid_Out & channel51_Kernel51_Valid_Out & channel52_Kernel51_Valid_Out & channel53_Kernel51_Valid_Out & channel54_Kernel51_Valid_Out & channel55_Kernel51_Valid_Out & channel56_Kernel51_Valid_Out & channel57_Kernel51_Valid_Out & channel58_Kernel51_Valid_Out & channel59_Kernel51_Valid_Out & channel60_Kernel51_Valid_Out & channel61_Kernel51_Valid_Out & channel62_Kernel51_Valid_Out & channel63_Kernel51_Valid_Out & channel64_Kernel51_Valid_Out;

	wire channel1_Kernel52_Valid_Out, channel2_Kernel52_Valid_Out, channel3_Kernel52_Valid_Out, channel4_Kernel52_Valid_Out, channel5_Kernel52_Valid_Out, channel6_Kernel52_Valid_Out, channel7_Kernel52_Valid_Out, channel8_Kernel52_Valid_Out, channel9_Kernel52_Valid_Out, channel10_Kernel52_Valid_Out, channel11_Kernel52_Valid_Out, channel12_Kernel52_Valid_Out, channel13_Kernel52_Valid_Out, channel14_Kernel52_Valid_Out, channel15_Kernel52_Valid_Out, channel16_Kernel52_Valid_Out, channel17_Kernel52_Valid_Out, channel18_Kernel52_Valid_Out, channel19_Kernel52_Valid_Out, channel20_Kernel52_Valid_Out, channel21_Kernel52_Valid_Out, channel22_Kernel52_Valid_Out, channel23_Kernel52_Valid_Out, channel24_Kernel52_Valid_Out, channel25_Kernel52_Valid_Out, channel26_Kernel52_Valid_Out, channel27_Kernel52_Valid_Out, channel28_Kernel52_Valid_Out, channel29_Kernel52_Valid_Out, channel30_Kernel52_Valid_Out, channel31_Kernel52_Valid_Out, channel32_Kernel52_Valid_Out, channel33_Kernel52_Valid_Out, channel34_Kernel52_Valid_Out, channel35_Kernel52_Valid_Out, channel36_Kernel52_Valid_Out, channel37_Kernel52_Valid_Out, channel38_Kernel52_Valid_Out, channel39_Kernel52_Valid_Out, channel40_Kernel52_Valid_Out, channel41_Kernel52_Valid_Out, channel42_Kernel52_Valid_Out, channel43_Kernel52_Valid_Out, channel44_Kernel52_Valid_Out, channel45_Kernel52_Valid_Out, channel46_Kernel52_Valid_Out, channel47_Kernel52_Valid_Out, channel48_Kernel52_Valid_Out, channel49_Kernel52_Valid_Out, channel50_Kernel52_Valid_Out, channel51_Kernel52_Valid_Out, channel52_Kernel52_Valid_Out, channel53_Kernel52_Valid_Out, channel54_Kernel52_Valid_Out, channel55_Kernel52_Valid_Out, channel56_Kernel52_Valid_Out, channel57_Kernel52_Valid_Out, channel58_Kernel52_Valid_Out, channel59_Kernel52_Valid_Out, channel60_Kernel52_Valid_Out, channel61_Kernel52_Valid_Out, channel62_Kernel52_Valid_Out, channel63_Kernel52_Valid_Out, channel64_Kernel52_Valid_Out;

	assign add_kernel52=channel1_Kernel52_Valid_Out & channel2_Kernel52_Valid_Out & channel3_Kernel52_Valid_Out & channel4_Kernel52_Valid_Out & channel5_Kernel52_Valid_Out & channel6_Kernel52_Valid_Out & channel7_Kernel52_Valid_Out & channel8_Kernel52_Valid_Out & channel9_Kernel52_Valid_Out & channel10_Kernel52_Valid_Out & channel11_Kernel52_Valid_Out & channel12_Kernel52_Valid_Out & channel13_Kernel52_Valid_Out & channel14_Kernel52_Valid_Out & channel15_Kernel52_Valid_Out & channel16_Kernel52_Valid_Out & channel17_Kernel52_Valid_Out & channel18_Kernel52_Valid_Out & channel19_Kernel52_Valid_Out & channel20_Kernel52_Valid_Out & channel21_Kernel52_Valid_Out & channel22_Kernel52_Valid_Out & channel23_Kernel52_Valid_Out & channel24_Kernel52_Valid_Out & channel25_Kernel52_Valid_Out & channel26_Kernel52_Valid_Out & channel27_Kernel52_Valid_Out & channel28_Kernel52_Valid_Out & channel29_Kernel52_Valid_Out & channel30_Kernel52_Valid_Out & channel31_Kernel52_Valid_Out & channel32_Kernel52_Valid_Out & channel33_Kernel52_Valid_Out & channel34_Kernel52_Valid_Out & channel35_Kernel52_Valid_Out & channel36_Kernel52_Valid_Out & channel37_Kernel52_Valid_Out & channel38_Kernel52_Valid_Out & channel39_Kernel52_Valid_Out & channel40_Kernel52_Valid_Out & channel41_Kernel52_Valid_Out & channel42_Kernel52_Valid_Out & channel43_Kernel52_Valid_Out & channel44_Kernel52_Valid_Out & channel45_Kernel52_Valid_Out & channel46_Kernel52_Valid_Out & channel47_Kernel52_Valid_Out & channel48_Kernel52_Valid_Out & channel49_Kernel52_Valid_Out & channel50_Kernel52_Valid_Out & channel51_Kernel52_Valid_Out & channel52_Kernel52_Valid_Out & channel53_Kernel52_Valid_Out & channel54_Kernel52_Valid_Out & channel55_Kernel52_Valid_Out & channel56_Kernel52_Valid_Out & channel57_Kernel52_Valid_Out & channel58_Kernel52_Valid_Out & channel59_Kernel52_Valid_Out & channel60_Kernel52_Valid_Out & channel61_Kernel52_Valid_Out & channel62_Kernel52_Valid_Out & channel63_Kernel52_Valid_Out & channel64_Kernel52_Valid_Out;

	wire channel1_Kernel53_Valid_Out, channel2_Kernel53_Valid_Out, channel3_Kernel53_Valid_Out, channel4_Kernel53_Valid_Out, channel5_Kernel53_Valid_Out, channel6_Kernel53_Valid_Out, channel7_Kernel53_Valid_Out, channel8_Kernel53_Valid_Out, channel9_Kernel53_Valid_Out, channel10_Kernel53_Valid_Out, channel11_Kernel53_Valid_Out, channel12_Kernel53_Valid_Out, channel13_Kernel53_Valid_Out, channel14_Kernel53_Valid_Out, channel15_Kernel53_Valid_Out, channel16_Kernel53_Valid_Out, channel17_Kernel53_Valid_Out, channel18_Kernel53_Valid_Out, channel19_Kernel53_Valid_Out, channel20_Kernel53_Valid_Out, channel21_Kernel53_Valid_Out, channel22_Kernel53_Valid_Out, channel23_Kernel53_Valid_Out, channel24_Kernel53_Valid_Out, channel25_Kernel53_Valid_Out, channel26_Kernel53_Valid_Out, channel27_Kernel53_Valid_Out, channel28_Kernel53_Valid_Out, channel29_Kernel53_Valid_Out, channel30_Kernel53_Valid_Out, channel31_Kernel53_Valid_Out, channel32_Kernel53_Valid_Out, channel33_Kernel53_Valid_Out, channel34_Kernel53_Valid_Out, channel35_Kernel53_Valid_Out, channel36_Kernel53_Valid_Out, channel37_Kernel53_Valid_Out, channel38_Kernel53_Valid_Out, channel39_Kernel53_Valid_Out, channel40_Kernel53_Valid_Out, channel41_Kernel53_Valid_Out, channel42_Kernel53_Valid_Out, channel43_Kernel53_Valid_Out, channel44_Kernel53_Valid_Out, channel45_Kernel53_Valid_Out, channel46_Kernel53_Valid_Out, channel47_Kernel53_Valid_Out, channel48_Kernel53_Valid_Out, channel49_Kernel53_Valid_Out, channel50_Kernel53_Valid_Out, channel51_Kernel53_Valid_Out, channel52_Kernel53_Valid_Out, channel53_Kernel53_Valid_Out, channel54_Kernel53_Valid_Out, channel55_Kernel53_Valid_Out, channel56_Kernel53_Valid_Out, channel57_Kernel53_Valid_Out, channel58_Kernel53_Valid_Out, channel59_Kernel53_Valid_Out, channel60_Kernel53_Valid_Out, channel61_Kernel53_Valid_Out, channel62_Kernel53_Valid_Out, channel63_Kernel53_Valid_Out, channel64_Kernel53_Valid_Out;

	assign add_kernel53=channel1_Kernel53_Valid_Out & channel2_Kernel53_Valid_Out & channel3_Kernel53_Valid_Out & channel4_Kernel53_Valid_Out & channel5_Kernel53_Valid_Out & channel6_Kernel53_Valid_Out & channel7_Kernel53_Valid_Out & channel8_Kernel53_Valid_Out & channel9_Kernel53_Valid_Out & channel10_Kernel53_Valid_Out & channel11_Kernel53_Valid_Out & channel12_Kernel53_Valid_Out & channel13_Kernel53_Valid_Out & channel14_Kernel53_Valid_Out & channel15_Kernel53_Valid_Out & channel16_Kernel53_Valid_Out & channel17_Kernel53_Valid_Out & channel18_Kernel53_Valid_Out & channel19_Kernel53_Valid_Out & channel20_Kernel53_Valid_Out & channel21_Kernel53_Valid_Out & channel22_Kernel53_Valid_Out & channel23_Kernel53_Valid_Out & channel24_Kernel53_Valid_Out & channel25_Kernel53_Valid_Out & channel26_Kernel53_Valid_Out & channel27_Kernel53_Valid_Out & channel28_Kernel53_Valid_Out & channel29_Kernel53_Valid_Out & channel30_Kernel53_Valid_Out & channel31_Kernel53_Valid_Out & channel32_Kernel53_Valid_Out & channel33_Kernel53_Valid_Out & channel34_Kernel53_Valid_Out & channel35_Kernel53_Valid_Out & channel36_Kernel53_Valid_Out & channel37_Kernel53_Valid_Out & channel38_Kernel53_Valid_Out & channel39_Kernel53_Valid_Out & channel40_Kernel53_Valid_Out & channel41_Kernel53_Valid_Out & channel42_Kernel53_Valid_Out & channel43_Kernel53_Valid_Out & channel44_Kernel53_Valid_Out & channel45_Kernel53_Valid_Out & channel46_Kernel53_Valid_Out & channel47_Kernel53_Valid_Out & channel48_Kernel53_Valid_Out & channel49_Kernel53_Valid_Out & channel50_Kernel53_Valid_Out & channel51_Kernel53_Valid_Out & channel52_Kernel53_Valid_Out & channel53_Kernel53_Valid_Out & channel54_Kernel53_Valid_Out & channel55_Kernel53_Valid_Out & channel56_Kernel53_Valid_Out & channel57_Kernel53_Valid_Out & channel58_Kernel53_Valid_Out & channel59_Kernel53_Valid_Out & channel60_Kernel53_Valid_Out & channel61_Kernel53_Valid_Out & channel62_Kernel53_Valid_Out & channel63_Kernel53_Valid_Out & channel64_Kernel53_Valid_Out;

	wire channel1_Kernel54_Valid_Out, channel2_Kernel54_Valid_Out, channel3_Kernel54_Valid_Out, channel4_Kernel54_Valid_Out, channel5_Kernel54_Valid_Out, channel6_Kernel54_Valid_Out, channel7_Kernel54_Valid_Out, channel8_Kernel54_Valid_Out, channel9_Kernel54_Valid_Out, channel10_Kernel54_Valid_Out, channel11_Kernel54_Valid_Out, channel12_Kernel54_Valid_Out, channel13_Kernel54_Valid_Out, channel14_Kernel54_Valid_Out, channel15_Kernel54_Valid_Out, channel16_Kernel54_Valid_Out, channel17_Kernel54_Valid_Out, channel18_Kernel54_Valid_Out, channel19_Kernel54_Valid_Out, channel20_Kernel54_Valid_Out, channel21_Kernel54_Valid_Out, channel22_Kernel54_Valid_Out, channel23_Kernel54_Valid_Out, channel24_Kernel54_Valid_Out, channel25_Kernel54_Valid_Out, channel26_Kernel54_Valid_Out, channel27_Kernel54_Valid_Out, channel28_Kernel54_Valid_Out, channel29_Kernel54_Valid_Out, channel30_Kernel54_Valid_Out, channel31_Kernel54_Valid_Out, channel32_Kernel54_Valid_Out, channel33_Kernel54_Valid_Out, channel34_Kernel54_Valid_Out, channel35_Kernel54_Valid_Out, channel36_Kernel54_Valid_Out, channel37_Kernel54_Valid_Out, channel38_Kernel54_Valid_Out, channel39_Kernel54_Valid_Out, channel40_Kernel54_Valid_Out, channel41_Kernel54_Valid_Out, channel42_Kernel54_Valid_Out, channel43_Kernel54_Valid_Out, channel44_Kernel54_Valid_Out, channel45_Kernel54_Valid_Out, channel46_Kernel54_Valid_Out, channel47_Kernel54_Valid_Out, channel48_Kernel54_Valid_Out, channel49_Kernel54_Valid_Out, channel50_Kernel54_Valid_Out, channel51_Kernel54_Valid_Out, channel52_Kernel54_Valid_Out, channel53_Kernel54_Valid_Out, channel54_Kernel54_Valid_Out, channel55_Kernel54_Valid_Out, channel56_Kernel54_Valid_Out, channel57_Kernel54_Valid_Out, channel58_Kernel54_Valid_Out, channel59_Kernel54_Valid_Out, channel60_Kernel54_Valid_Out, channel61_Kernel54_Valid_Out, channel62_Kernel54_Valid_Out, channel63_Kernel54_Valid_Out, channel64_Kernel54_Valid_Out;

	assign add_kernel54=channel1_Kernel54_Valid_Out & channel2_Kernel54_Valid_Out & channel3_Kernel54_Valid_Out & channel4_Kernel54_Valid_Out & channel5_Kernel54_Valid_Out & channel6_Kernel54_Valid_Out & channel7_Kernel54_Valid_Out & channel8_Kernel54_Valid_Out & channel9_Kernel54_Valid_Out & channel10_Kernel54_Valid_Out & channel11_Kernel54_Valid_Out & channel12_Kernel54_Valid_Out & channel13_Kernel54_Valid_Out & channel14_Kernel54_Valid_Out & channel15_Kernel54_Valid_Out & channel16_Kernel54_Valid_Out & channel17_Kernel54_Valid_Out & channel18_Kernel54_Valid_Out & channel19_Kernel54_Valid_Out & channel20_Kernel54_Valid_Out & channel21_Kernel54_Valid_Out & channel22_Kernel54_Valid_Out & channel23_Kernel54_Valid_Out & channel24_Kernel54_Valid_Out & channel25_Kernel54_Valid_Out & channel26_Kernel54_Valid_Out & channel27_Kernel54_Valid_Out & channel28_Kernel54_Valid_Out & channel29_Kernel54_Valid_Out & channel30_Kernel54_Valid_Out & channel31_Kernel54_Valid_Out & channel32_Kernel54_Valid_Out & channel33_Kernel54_Valid_Out & channel34_Kernel54_Valid_Out & channel35_Kernel54_Valid_Out & channel36_Kernel54_Valid_Out & channel37_Kernel54_Valid_Out & channel38_Kernel54_Valid_Out & channel39_Kernel54_Valid_Out & channel40_Kernel54_Valid_Out & channel41_Kernel54_Valid_Out & channel42_Kernel54_Valid_Out & channel43_Kernel54_Valid_Out & channel44_Kernel54_Valid_Out & channel45_Kernel54_Valid_Out & channel46_Kernel54_Valid_Out & channel47_Kernel54_Valid_Out & channel48_Kernel54_Valid_Out & channel49_Kernel54_Valid_Out & channel50_Kernel54_Valid_Out & channel51_Kernel54_Valid_Out & channel52_Kernel54_Valid_Out & channel53_Kernel54_Valid_Out & channel54_Kernel54_Valid_Out & channel55_Kernel54_Valid_Out & channel56_Kernel54_Valid_Out & channel57_Kernel54_Valid_Out & channel58_Kernel54_Valid_Out & channel59_Kernel54_Valid_Out & channel60_Kernel54_Valid_Out & channel61_Kernel54_Valid_Out & channel62_Kernel54_Valid_Out & channel63_Kernel54_Valid_Out & channel64_Kernel54_Valid_Out;

	wire channel1_Kernel55_Valid_Out, channel2_Kernel55_Valid_Out, channel3_Kernel55_Valid_Out, channel4_Kernel55_Valid_Out, channel5_Kernel55_Valid_Out, channel6_Kernel55_Valid_Out, channel7_Kernel55_Valid_Out, channel8_Kernel55_Valid_Out, channel9_Kernel55_Valid_Out, channel10_Kernel55_Valid_Out, channel11_Kernel55_Valid_Out, channel12_Kernel55_Valid_Out, channel13_Kernel55_Valid_Out, channel14_Kernel55_Valid_Out, channel15_Kernel55_Valid_Out, channel16_Kernel55_Valid_Out, channel17_Kernel55_Valid_Out, channel18_Kernel55_Valid_Out, channel19_Kernel55_Valid_Out, channel20_Kernel55_Valid_Out, channel21_Kernel55_Valid_Out, channel22_Kernel55_Valid_Out, channel23_Kernel55_Valid_Out, channel24_Kernel55_Valid_Out, channel25_Kernel55_Valid_Out, channel26_Kernel55_Valid_Out, channel27_Kernel55_Valid_Out, channel28_Kernel55_Valid_Out, channel29_Kernel55_Valid_Out, channel30_Kernel55_Valid_Out, channel31_Kernel55_Valid_Out, channel32_Kernel55_Valid_Out, channel33_Kernel55_Valid_Out, channel34_Kernel55_Valid_Out, channel35_Kernel55_Valid_Out, channel36_Kernel55_Valid_Out, channel37_Kernel55_Valid_Out, channel38_Kernel55_Valid_Out, channel39_Kernel55_Valid_Out, channel40_Kernel55_Valid_Out, channel41_Kernel55_Valid_Out, channel42_Kernel55_Valid_Out, channel43_Kernel55_Valid_Out, channel44_Kernel55_Valid_Out, channel45_Kernel55_Valid_Out, channel46_Kernel55_Valid_Out, channel47_Kernel55_Valid_Out, channel48_Kernel55_Valid_Out, channel49_Kernel55_Valid_Out, channel50_Kernel55_Valid_Out, channel51_Kernel55_Valid_Out, channel52_Kernel55_Valid_Out, channel53_Kernel55_Valid_Out, channel54_Kernel55_Valid_Out, channel55_Kernel55_Valid_Out, channel56_Kernel55_Valid_Out, channel57_Kernel55_Valid_Out, channel58_Kernel55_Valid_Out, channel59_Kernel55_Valid_Out, channel60_Kernel55_Valid_Out, channel61_Kernel55_Valid_Out, channel62_Kernel55_Valid_Out, channel63_Kernel55_Valid_Out, channel64_Kernel55_Valid_Out;

	assign add_kernel55=channel1_Kernel55_Valid_Out & channel2_Kernel55_Valid_Out & channel3_Kernel55_Valid_Out & channel4_Kernel55_Valid_Out & channel5_Kernel55_Valid_Out & channel6_Kernel55_Valid_Out & channel7_Kernel55_Valid_Out & channel8_Kernel55_Valid_Out & channel9_Kernel55_Valid_Out & channel10_Kernel55_Valid_Out & channel11_Kernel55_Valid_Out & channel12_Kernel55_Valid_Out & channel13_Kernel55_Valid_Out & channel14_Kernel55_Valid_Out & channel15_Kernel55_Valid_Out & channel16_Kernel55_Valid_Out & channel17_Kernel55_Valid_Out & channel18_Kernel55_Valid_Out & channel19_Kernel55_Valid_Out & channel20_Kernel55_Valid_Out & channel21_Kernel55_Valid_Out & channel22_Kernel55_Valid_Out & channel23_Kernel55_Valid_Out & channel24_Kernel55_Valid_Out & channel25_Kernel55_Valid_Out & channel26_Kernel55_Valid_Out & channel27_Kernel55_Valid_Out & channel28_Kernel55_Valid_Out & channel29_Kernel55_Valid_Out & channel30_Kernel55_Valid_Out & channel31_Kernel55_Valid_Out & channel32_Kernel55_Valid_Out & channel33_Kernel55_Valid_Out & channel34_Kernel55_Valid_Out & channel35_Kernel55_Valid_Out & channel36_Kernel55_Valid_Out & channel37_Kernel55_Valid_Out & channel38_Kernel55_Valid_Out & channel39_Kernel55_Valid_Out & channel40_Kernel55_Valid_Out & channel41_Kernel55_Valid_Out & channel42_Kernel55_Valid_Out & channel43_Kernel55_Valid_Out & channel44_Kernel55_Valid_Out & channel45_Kernel55_Valid_Out & channel46_Kernel55_Valid_Out & channel47_Kernel55_Valid_Out & channel48_Kernel55_Valid_Out & channel49_Kernel55_Valid_Out & channel50_Kernel55_Valid_Out & channel51_Kernel55_Valid_Out & channel52_Kernel55_Valid_Out & channel53_Kernel55_Valid_Out & channel54_Kernel55_Valid_Out & channel55_Kernel55_Valid_Out & channel56_Kernel55_Valid_Out & channel57_Kernel55_Valid_Out & channel58_Kernel55_Valid_Out & channel59_Kernel55_Valid_Out & channel60_Kernel55_Valid_Out & channel61_Kernel55_Valid_Out & channel62_Kernel55_Valid_Out & channel63_Kernel55_Valid_Out & channel64_Kernel55_Valid_Out;

	wire channel1_Kernel56_Valid_Out, channel2_Kernel56_Valid_Out, channel3_Kernel56_Valid_Out, channel4_Kernel56_Valid_Out, channel5_Kernel56_Valid_Out, channel6_Kernel56_Valid_Out, channel7_Kernel56_Valid_Out, channel8_Kernel56_Valid_Out, channel9_Kernel56_Valid_Out, channel10_Kernel56_Valid_Out, channel11_Kernel56_Valid_Out, channel12_Kernel56_Valid_Out, channel13_Kernel56_Valid_Out, channel14_Kernel56_Valid_Out, channel15_Kernel56_Valid_Out, channel16_Kernel56_Valid_Out, channel17_Kernel56_Valid_Out, channel18_Kernel56_Valid_Out, channel19_Kernel56_Valid_Out, channel20_Kernel56_Valid_Out, channel21_Kernel56_Valid_Out, channel22_Kernel56_Valid_Out, channel23_Kernel56_Valid_Out, channel24_Kernel56_Valid_Out, channel25_Kernel56_Valid_Out, channel26_Kernel56_Valid_Out, channel27_Kernel56_Valid_Out, channel28_Kernel56_Valid_Out, channel29_Kernel56_Valid_Out, channel30_Kernel56_Valid_Out, channel31_Kernel56_Valid_Out, channel32_Kernel56_Valid_Out, channel33_Kernel56_Valid_Out, channel34_Kernel56_Valid_Out, channel35_Kernel56_Valid_Out, channel36_Kernel56_Valid_Out, channel37_Kernel56_Valid_Out, channel38_Kernel56_Valid_Out, channel39_Kernel56_Valid_Out, channel40_Kernel56_Valid_Out, channel41_Kernel56_Valid_Out, channel42_Kernel56_Valid_Out, channel43_Kernel56_Valid_Out, channel44_Kernel56_Valid_Out, channel45_Kernel56_Valid_Out, channel46_Kernel56_Valid_Out, channel47_Kernel56_Valid_Out, channel48_Kernel56_Valid_Out, channel49_Kernel56_Valid_Out, channel50_Kernel56_Valid_Out, channel51_Kernel56_Valid_Out, channel52_Kernel56_Valid_Out, channel53_Kernel56_Valid_Out, channel54_Kernel56_Valid_Out, channel55_Kernel56_Valid_Out, channel56_Kernel56_Valid_Out, channel57_Kernel56_Valid_Out, channel58_Kernel56_Valid_Out, channel59_Kernel56_Valid_Out, channel60_Kernel56_Valid_Out, channel61_Kernel56_Valid_Out, channel62_Kernel56_Valid_Out, channel63_Kernel56_Valid_Out, channel64_Kernel56_Valid_Out;

	assign add_kernel56=channel1_Kernel56_Valid_Out & channel2_Kernel56_Valid_Out & channel3_Kernel56_Valid_Out & channel4_Kernel56_Valid_Out & channel5_Kernel56_Valid_Out & channel6_Kernel56_Valid_Out & channel7_Kernel56_Valid_Out & channel8_Kernel56_Valid_Out & channel9_Kernel56_Valid_Out & channel10_Kernel56_Valid_Out & channel11_Kernel56_Valid_Out & channel12_Kernel56_Valid_Out & channel13_Kernel56_Valid_Out & channel14_Kernel56_Valid_Out & channel15_Kernel56_Valid_Out & channel16_Kernel56_Valid_Out & channel17_Kernel56_Valid_Out & channel18_Kernel56_Valid_Out & channel19_Kernel56_Valid_Out & channel20_Kernel56_Valid_Out & channel21_Kernel56_Valid_Out & channel22_Kernel56_Valid_Out & channel23_Kernel56_Valid_Out & channel24_Kernel56_Valid_Out & channel25_Kernel56_Valid_Out & channel26_Kernel56_Valid_Out & channel27_Kernel56_Valid_Out & channel28_Kernel56_Valid_Out & channel29_Kernel56_Valid_Out & channel30_Kernel56_Valid_Out & channel31_Kernel56_Valid_Out & channel32_Kernel56_Valid_Out & channel33_Kernel56_Valid_Out & channel34_Kernel56_Valid_Out & channel35_Kernel56_Valid_Out & channel36_Kernel56_Valid_Out & channel37_Kernel56_Valid_Out & channel38_Kernel56_Valid_Out & channel39_Kernel56_Valid_Out & channel40_Kernel56_Valid_Out & channel41_Kernel56_Valid_Out & channel42_Kernel56_Valid_Out & channel43_Kernel56_Valid_Out & channel44_Kernel56_Valid_Out & channel45_Kernel56_Valid_Out & channel46_Kernel56_Valid_Out & channel47_Kernel56_Valid_Out & channel48_Kernel56_Valid_Out & channel49_Kernel56_Valid_Out & channel50_Kernel56_Valid_Out & channel51_Kernel56_Valid_Out & channel52_Kernel56_Valid_Out & channel53_Kernel56_Valid_Out & channel54_Kernel56_Valid_Out & channel55_Kernel56_Valid_Out & channel56_Kernel56_Valid_Out & channel57_Kernel56_Valid_Out & channel58_Kernel56_Valid_Out & channel59_Kernel56_Valid_Out & channel60_Kernel56_Valid_Out & channel61_Kernel56_Valid_Out & channel62_Kernel56_Valid_Out & channel63_Kernel56_Valid_Out & channel64_Kernel56_Valid_Out;

	wire channel1_Kernel57_Valid_Out, channel2_Kernel57_Valid_Out, channel3_Kernel57_Valid_Out, channel4_Kernel57_Valid_Out, channel5_Kernel57_Valid_Out, channel6_Kernel57_Valid_Out, channel7_Kernel57_Valid_Out, channel8_Kernel57_Valid_Out, channel9_Kernel57_Valid_Out, channel10_Kernel57_Valid_Out, channel11_Kernel57_Valid_Out, channel12_Kernel57_Valid_Out, channel13_Kernel57_Valid_Out, channel14_Kernel57_Valid_Out, channel15_Kernel57_Valid_Out, channel16_Kernel57_Valid_Out, channel17_Kernel57_Valid_Out, channel18_Kernel57_Valid_Out, channel19_Kernel57_Valid_Out, channel20_Kernel57_Valid_Out, channel21_Kernel57_Valid_Out, channel22_Kernel57_Valid_Out, channel23_Kernel57_Valid_Out, channel24_Kernel57_Valid_Out, channel25_Kernel57_Valid_Out, channel26_Kernel57_Valid_Out, channel27_Kernel57_Valid_Out, channel28_Kernel57_Valid_Out, channel29_Kernel57_Valid_Out, channel30_Kernel57_Valid_Out, channel31_Kernel57_Valid_Out, channel32_Kernel57_Valid_Out, channel33_Kernel57_Valid_Out, channel34_Kernel57_Valid_Out, channel35_Kernel57_Valid_Out, channel36_Kernel57_Valid_Out, channel37_Kernel57_Valid_Out, channel38_Kernel57_Valid_Out, channel39_Kernel57_Valid_Out, channel40_Kernel57_Valid_Out, channel41_Kernel57_Valid_Out, channel42_Kernel57_Valid_Out, channel43_Kernel57_Valid_Out, channel44_Kernel57_Valid_Out, channel45_Kernel57_Valid_Out, channel46_Kernel57_Valid_Out, channel47_Kernel57_Valid_Out, channel48_Kernel57_Valid_Out, channel49_Kernel57_Valid_Out, channel50_Kernel57_Valid_Out, channel51_Kernel57_Valid_Out, channel52_Kernel57_Valid_Out, channel53_Kernel57_Valid_Out, channel54_Kernel57_Valid_Out, channel55_Kernel57_Valid_Out, channel56_Kernel57_Valid_Out, channel57_Kernel57_Valid_Out, channel58_Kernel57_Valid_Out, channel59_Kernel57_Valid_Out, channel60_Kernel57_Valid_Out, channel61_Kernel57_Valid_Out, channel62_Kernel57_Valid_Out, channel63_Kernel57_Valid_Out, channel64_Kernel57_Valid_Out;

	assign add_kernel57=channel1_Kernel57_Valid_Out & channel2_Kernel57_Valid_Out & channel3_Kernel57_Valid_Out & channel4_Kernel57_Valid_Out & channel5_Kernel57_Valid_Out & channel6_Kernel57_Valid_Out & channel7_Kernel57_Valid_Out & channel8_Kernel57_Valid_Out & channel9_Kernel57_Valid_Out & channel10_Kernel57_Valid_Out & channel11_Kernel57_Valid_Out & channel12_Kernel57_Valid_Out & channel13_Kernel57_Valid_Out & channel14_Kernel57_Valid_Out & channel15_Kernel57_Valid_Out & channel16_Kernel57_Valid_Out & channel17_Kernel57_Valid_Out & channel18_Kernel57_Valid_Out & channel19_Kernel57_Valid_Out & channel20_Kernel57_Valid_Out & channel21_Kernel57_Valid_Out & channel22_Kernel57_Valid_Out & channel23_Kernel57_Valid_Out & channel24_Kernel57_Valid_Out & channel25_Kernel57_Valid_Out & channel26_Kernel57_Valid_Out & channel27_Kernel57_Valid_Out & channel28_Kernel57_Valid_Out & channel29_Kernel57_Valid_Out & channel30_Kernel57_Valid_Out & channel31_Kernel57_Valid_Out & channel32_Kernel57_Valid_Out & channel33_Kernel57_Valid_Out & channel34_Kernel57_Valid_Out & channel35_Kernel57_Valid_Out & channel36_Kernel57_Valid_Out & channel37_Kernel57_Valid_Out & channel38_Kernel57_Valid_Out & channel39_Kernel57_Valid_Out & channel40_Kernel57_Valid_Out & channel41_Kernel57_Valid_Out & channel42_Kernel57_Valid_Out & channel43_Kernel57_Valid_Out & channel44_Kernel57_Valid_Out & channel45_Kernel57_Valid_Out & channel46_Kernel57_Valid_Out & channel47_Kernel57_Valid_Out & channel48_Kernel57_Valid_Out & channel49_Kernel57_Valid_Out & channel50_Kernel57_Valid_Out & channel51_Kernel57_Valid_Out & channel52_Kernel57_Valid_Out & channel53_Kernel57_Valid_Out & channel54_Kernel57_Valid_Out & channel55_Kernel57_Valid_Out & channel56_Kernel57_Valid_Out & channel57_Kernel57_Valid_Out & channel58_Kernel57_Valid_Out & channel59_Kernel57_Valid_Out & channel60_Kernel57_Valid_Out & channel61_Kernel57_Valid_Out & channel62_Kernel57_Valid_Out & channel63_Kernel57_Valid_Out & channel64_Kernel57_Valid_Out;

	wire channel1_Kernel58_Valid_Out, channel2_Kernel58_Valid_Out, channel3_Kernel58_Valid_Out, channel4_Kernel58_Valid_Out, channel5_Kernel58_Valid_Out, channel6_Kernel58_Valid_Out, channel7_Kernel58_Valid_Out, channel8_Kernel58_Valid_Out, channel9_Kernel58_Valid_Out, channel10_Kernel58_Valid_Out, channel11_Kernel58_Valid_Out, channel12_Kernel58_Valid_Out, channel13_Kernel58_Valid_Out, channel14_Kernel58_Valid_Out, channel15_Kernel58_Valid_Out, channel16_Kernel58_Valid_Out, channel17_Kernel58_Valid_Out, channel18_Kernel58_Valid_Out, channel19_Kernel58_Valid_Out, channel20_Kernel58_Valid_Out, channel21_Kernel58_Valid_Out, channel22_Kernel58_Valid_Out, channel23_Kernel58_Valid_Out, channel24_Kernel58_Valid_Out, channel25_Kernel58_Valid_Out, channel26_Kernel58_Valid_Out, channel27_Kernel58_Valid_Out, channel28_Kernel58_Valid_Out, channel29_Kernel58_Valid_Out, channel30_Kernel58_Valid_Out, channel31_Kernel58_Valid_Out, channel32_Kernel58_Valid_Out, channel33_Kernel58_Valid_Out, channel34_Kernel58_Valid_Out, channel35_Kernel58_Valid_Out, channel36_Kernel58_Valid_Out, channel37_Kernel58_Valid_Out, channel38_Kernel58_Valid_Out, channel39_Kernel58_Valid_Out, channel40_Kernel58_Valid_Out, channel41_Kernel58_Valid_Out, channel42_Kernel58_Valid_Out, channel43_Kernel58_Valid_Out, channel44_Kernel58_Valid_Out, channel45_Kernel58_Valid_Out, channel46_Kernel58_Valid_Out, channel47_Kernel58_Valid_Out, channel48_Kernel58_Valid_Out, channel49_Kernel58_Valid_Out, channel50_Kernel58_Valid_Out, channel51_Kernel58_Valid_Out, channel52_Kernel58_Valid_Out, channel53_Kernel58_Valid_Out, channel54_Kernel58_Valid_Out, channel55_Kernel58_Valid_Out, channel56_Kernel58_Valid_Out, channel57_Kernel58_Valid_Out, channel58_Kernel58_Valid_Out, channel59_Kernel58_Valid_Out, channel60_Kernel58_Valid_Out, channel61_Kernel58_Valid_Out, channel62_Kernel58_Valid_Out, channel63_Kernel58_Valid_Out, channel64_Kernel58_Valid_Out;

	assign add_kernel58=channel1_Kernel58_Valid_Out & channel2_Kernel58_Valid_Out & channel3_Kernel58_Valid_Out & channel4_Kernel58_Valid_Out & channel5_Kernel58_Valid_Out & channel6_Kernel58_Valid_Out & channel7_Kernel58_Valid_Out & channel8_Kernel58_Valid_Out & channel9_Kernel58_Valid_Out & channel10_Kernel58_Valid_Out & channel11_Kernel58_Valid_Out & channel12_Kernel58_Valid_Out & channel13_Kernel58_Valid_Out & channel14_Kernel58_Valid_Out & channel15_Kernel58_Valid_Out & channel16_Kernel58_Valid_Out & channel17_Kernel58_Valid_Out & channel18_Kernel58_Valid_Out & channel19_Kernel58_Valid_Out & channel20_Kernel58_Valid_Out & channel21_Kernel58_Valid_Out & channel22_Kernel58_Valid_Out & channel23_Kernel58_Valid_Out & channel24_Kernel58_Valid_Out & channel25_Kernel58_Valid_Out & channel26_Kernel58_Valid_Out & channel27_Kernel58_Valid_Out & channel28_Kernel58_Valid_Out & channel29_Kernel58_Valid_Out & channel30_Kernel58_Valid_Out & channel31_Kernel58_Valid_Out & channel32_Kernel58_Valid_Out & channel33_Kernel58_Valid_Out & channel34_Kernel58_Valid_Out & channel35_Kernel58_Valid_Out & channel36_Kernel58_Valid_Out & channel37_Kernel58_Valid_Out & channel38_Kernel58_Valid_Out & channel39_Kernel58_Valid_Out & channel40_Kernel58_Valid_Out & channel41_Kernel58_Valid_Out & channel42_Kernel58_Valid_Out & channel43_Kernel58_Valid_Out & channel44_Kernel58_Valid_Out & channel45_Kernel58_Valid_Out & channel46_Kernel58_Valid_Out & channel47_Kernel58_Valid_Out & channel48_Kernel58_Valid_Out & channel49_Kernel58_Valid_Out & channel50_Kernel58_Valid_Out & channel51_Kernel58_Valid_Out & channel52_Kernel58_Valid_Out & channel53_Kernel58_Valid_Out & channel54_Kernel58_Valid_Out & channel55_Kernel58_Valid_Out & channel56_Kernel58_Valid_Out & channel57_Kernel58_Valid_Out & channel58_Kernel58_Valid_Out & channel59_Kernel58_Valid_Out & channel60_Kernel58_Valid_Out & channel61_Kernel58_Valid_Out & channel62_Kernel58_Valid_Out & channel63_Kernel58_Valid_Out & channel64_Kernel58_Valid_Out;

	wire channel1_Kernel59_Valid_Out, channel2_Kernel59_Valid_Out, channel3_Kernel59_Valid_Out, channel4_Kernel59_Valid_Out, channel5_Kernel59_Valid_Out, channel6_Kernel59_Valid_Out, channel7_Kernel59_Valid_Out, channel8_Kernel59_Valid_Out, channel9_Kernel59_Valid_Out, channel10_Kernel59_Valid_Out, channel11_Kernel59_Valid_Out, channel12_Kernel59_Valid_Out, channel13_Kernel59_Valid_Out, channel14_Kernel59_Valid_Out, channel15_Kernel59_Valid_Out, channel16_Kernel59_Valid_Out, channel17_Kernel59_Valid_Out, channel18_Kernel59_Valid_Out, channel19_Kernel59_Valid_Out, channel20_Kernel59_Valid_Out, channel21_Kernel59_Valid_Out, channel22_Kernel59_Valid_Out, channel23_Kernel59_Valid_Out, channel24_Kernel59_Valid_Out, channel25_Kernel59_Valid_Out, channel26_Kernel59_Valid_Out, channel27_Kernel59_Valid_Out, channel28_Kernel59_Valid_Out, channel29_Kernel59_Valid_Out, channel30_Kernel59_Valid_Out, channel31_Kernel59_Valid_Out, channel32_Kernel59_Valid_Out, channel33_Kernel59_Valid_Out, channel34_Kernel59_Valid_Out, channel35_Kernel59_Valid_Out, channel36_Kernel59_Valid_Out, channel37_Kernel59_Valid_Out, channel38_Kernel59_Valid_Out, channel39_Kernel59_Valid_Out, channel40_Kernel59_Valid_Out, channel41_Kernel59_Valid_Out, channel42_Kernel59_Valid_Out, channel43_Kernel59_Valid_Out, channel44_Kernel59_Valid_Out, channel45_Kernel59_Valid_Out, channel46_Kernel59_Valid_Out, channel47_Kernel59_Valid_Out, channel48_Kernel59_Valid_Out, channel49_Kernel59_Valid_Out, channel50_Kernel59_Valid_Out, channel51_Kernel59_Valid_Out, channel52_Kernel59_Valid_Out, channel53_Kernel59_Valid_Out, channel54_Kernel59_Valid_Out, channel55_Kernel59_Valid_Out, channel56_Kernel59_Valid_Out, channel57_Kernel59_Valid_Out, channel58_Kernel59_Valid_Out, channel59_Kernel59_Valid_Out, channel60_Kernel59_Valid_Out, channel61_Kernel59_Valid_Out, channel62_Kernel59_Valid_Out, channel63_Kernel59_Valid_Out, channel64_Kernel59_Valid_Out;

	assign add_kernel59=channel1_Kernel59_Valid_Out & channel2_Kernel59_Valid_Out & channel3_Kernel59_Valid_Out & channel4_Kernel59_Valid_Out & channel5_Kernel59_Valid_Out & channel6_Kernel59_Valid_Out & channel7_Kernel59_Valid_Out & channel8_Kernel59_Valid_Out & channel9_Kernel59_Valid_Out & channel10_Kernel59_Valid_Out & channel11_Kernel59_Valid_Out & channel12_Kernel59_Valid_Out & channel13_Kernel59_Valid_Out & channel14_Kernel59_Valid_Out & channel15_Kernel59_Valid_Out & channel16_Kernel59_Valid_Out & channel17_Kernel59_Valid_Out & channel18_Kernel59_Valid_Out & channel19_Kernel59_Valid_Out & channel20_Kernel59_Valid_Out & channel21_Kernel59_Valid_Out & channel22_Kernel59_Valid_Out & channel23_Kernel59_Valid_Out & channel24_Kernel59_Valid_Out & channel25_Kernel59_Valid_Out & channel26_Kernel59_Valid_Out & channel27_Kernel59_Valid_Out & channel28_Kernel59_Valid_Out & channel29_Kernel59_Valid_Out & channel30_Kernel59_Valid_Out & channel31_Kernel59_Valid_Out & channel32_Kernel59_Valid_Out & channel33_Kernel59_Valid_Out & channel34_Kernel59_Valid_Out & channel35_Kernel59_Valid_Out & channel36_Kernel59_Valid_Out & channel37_Kernel59_Valid_Out & channel38_Kernel59_Valid_Out & channel39_Kernel59_Valid_Out & channel40_Kernel59_Valid_Out & channel41_Kernel59_Valid_Out & channel42_Kernel59_Valid_Out & channel43_Kernel59_Valid_Out & channel44_Kernel59_Valid_Out & channel45_Kernel59_Valid_Out & channel46_Kernel59_Valid_Out & channel47_Kernel59_Valid_Out & channel48_Kernel59_Valid_Out & channel49_Kernel59_Valid_Out & channel50_Kernel59_Valid_Out & channel51_Kernel59_Valid_Out & channel52_Kernel59_Valid_Out & channel53_Kernel59_Valid_Out & channel54_Kernel59_Valid_Out & channel55_Kernel59_Valid_Out & channel56_Kernel59_Valid_Out & channel57_Kernel59_Valid_Out & channel58_Kernel59_Valid_Out & channel59_Kernel59_Valid_Out & channel60_Kernel59_Valid_Out & channel61_Kernel59_Valid_Out & channel62_Kernel59_Valid_Out & channel63_Kernel59_Valid_Out & channel64_Kernel59_Valid_Out;

	wire channel1_Kernel60_Valid_Out, channel2_Kernel60_Valid_Out, channel3_Kernel60_Valid_Out, channel4_Kernel60_Valid_Out, channel5_Kernel60_Valid_Out, channel6_Kernel60_Valid_Out, channel7_Kernel60_Valid_Out, channel8_Kernel60_Valid_Out, channel9_Kernel60_Valid_Out, channel10_Kernel60_Valid_Out, channel11_Kernel60_Valid_Out, channel12_Kernel60_Valid_Out, channel13_Kernel60_Valid_Out, channel14_Kernel60_Valid_Out, channel15_Kernel60_Valid_Out, channel16_Kernel60_Valid_Out, channel17_Kernel60_Valid_Out, channel18_Kernel60_Valid_Out, channel19_Kernel60_Valid_Out, channel20_Kernel60_Valid_Out, channel21_Kernel60_Valid_Out, channel22_Kernel60_Valid_Out, channel23_Kernel60_Valid_Out, channel24_Kernel60_Valid_Out, channel25_Kernel60_Valid_Out, channel26_Kernel60_Valid_Out, channel27_Kernel60_Valid_Out, channel28_Kernel60_Valid_Out, channel29_Kernel60_Valid_Out, channel30_Kernel60_Valid_Out, channel31_Kernel60_Valid_Out, channel32_Kernel60_Valid_Out, channel33_Kernel60_Valid_Out, channel34_Kernel60_Valid_Out, channel35_Kernel60_Valid_Out, channel36_Kernel60_Valid_Out, channel37_Kernel60_Valid_Out, channel38_Kernel60_Valid_Out, channel39_Kernel60_Valid_Out, channel40_Kernel60_Valid_Out, channel41_Kernel60_Valid_Out, channel42_Kernel60_Valid_Out, channel43_Kernel60_Valid_Out, channel44_Kernel60_Valid_Out, channel45_Kernel60_Valid_Out, channel46_Kernel60_Valid_Out, channel47_Kernel60_Valid_Out, channel48_Kernel60_Valid_Out, channel49_Kernel60_Valid_Out, channel50_Kernel60_Valid_Out, channel51_Kernel60_Valid_Out, channel52_Kernel60_Valid_Out, channel53_Kernel60_Valid_Out, channel54_Kernel60_Valid_Out, channel55_Kernel60_Valid_Out, channel56_Kernel60_Valid_Out, channel57_Kernel60_Valid_Out, channel58_Kernel60_Valid_Out, channel59_Kernel60_Valid_Out, channel60_Kernel60_Valid_Out, channel61_Kernel60_Valid_Out, channel62_Kernel60_Valid_Out, channel63_Kernel60_Valid_Out, channel64_Kernel60_Valid_Out;

	assign add_kernel60=channel1_Kernel60_Valid_Out & channel2_Kernel60_Valid_Out & channel3_Kernel60_Valid_Out & channel4_Kernel60_Valid_Out & channel5_Kernel60_Valid_Out & channel6_Kernel60_Valid_Out & channel7_Kernel60_Valid_Out & channel8_Kernel60_Valid_Out & channel9_Kernel60_Valid_Out & channel10_Kernel60_Valid_Out & channel11_Kernel60_Valid_Out & channel12_Kernel60_Valid_Out & channel13_Kernel60_Valid_Out & channel14_Kernel60_Valid_Out & channel15_Kernel60_Valid_Out & channel16_Kernel60_Valid_Out & channel17_Kernel60_Valid_Out & channel18_Kernel60_Valid_Out & channel19_Kernel60_Valid_Out & channel20_Kernel60_Valid_Out & channel21_Kernel60_Valid_Out & channel22_Kernel60_Valid_Out & channel23_Kernel60_Valid_Out & channel24_Kernel60_Valid_Out & channel25_Kernel60_Valid_Out & channel26_Kernel60_Valid_Out & channel27_Kernel60_Valid_Out & channel28_Kernel60_Valid_Out & channel29_Kernel60_Valid_Out & channel30_Kernel60_Valid_Out & channel31_Kernel60_Valid_Out & channel32_Kernel60_Valid_Out & channel33_Kernel60_Valid_Out & channel34_Kernel60_Valid_Out & channel35_Kernel60_Valid_Out & channel36_Kernel60_Valid_Out & channel37_Kernel60_Valid_Out & channel38_Kernel60_Valid_Out & channel39_Kernel60_Valid_Out & channel40_Kernel60_Valid_Out & channel41_Kernel60_Valid_Out & channel42_Kernel60_Valid_Out & channel43_Kernel60_Valid_Out & channel44_Kernel60_Valid_Out & channel45_Kernel60_Valid_Out & channel46_Kernel60_Valid_Out & channel47_Kernel60_Valid_Out & channel48_Kernel60_Valid_Out & channel49_Kernel60_Valid_Out & channel50_Kernel60_Valid_Out & channel51_Kernel60_Valid_Out & channel52_Kernel60_Valid_Out & channel53_Kernel60_Valid_Out & channel54_Kernel60_Valid_Out & channel55_Kernel60_Valid_Out & channel56_Kernel60_Valid_Out & channel57_Kernel60_Valid_Out & channel58_Kernel60_Valid_Out & channel59_Kernel60_Valid_Out & channel60_Kernel60_Valid_Out & channel61_Kernel60_Valid_Out & channel62_Kernel60_Valid_Out & channel63_Kernel60_Valid_Out & channel64_Kernel60_Valid_Out;

	wire channel1_Kernel61_Valid_Out, channel2_Kernel61_Valid_Out, channel3_Kernel61_Valid_Out, channel4_Kernel61_Valid_Out, channel5_Kernel61_Valid_Out, channel6_Kernel61_Valid_Out, channel7_Kernel61_Valid_Out, channel8_Kernel61_Valid_Out, channel9_Kernel61_Valid_Out, channel10_Kernel61_Valid_Out, channel11_Kernel61_Valid_Out, channel12_Kernel61_Valid_Out, channel13_Kernel61_Valid_Out, channel14_Kernel61_Valid_Out, channel15_Kernel61_Valid_Out, channel16_Kernel61_Valid_Out, channel17_Kernel61_Valid_Out, channel18_Kernel61_Valid_Out, channel19_Kernel61_Valid_Out, channel20_Kernel61_Valid_Out, channel21_Kernel61_Valid_Out, channel22_Kernel61_Valid_Out, channel23_Kernel61_Valid_Out, channel24_Kernel61_Valid_Out, channel25_Kernel61_Valid_Out, channel26_Kernel61_Valid_Out, channel27_Kernel61_Valid_Out, channel28_Kernel61_Valid_Out, channel29_Kernel61_Valid_Out, channel30_Kernel61_Valid_Out, channel31_Kernel61_Valid_Out, channel32_Kernel61_Valid_Out, channel33_Kernel61_Valid_Out, channel34_Kernel61_Valid_Out, channel35_Kernel61_Valid_Out, channel36_Kernel61_Valid_Out, channel37_Kernel61_Valid_Out, channel38_Kernel61_Valid_Out, channel39_Kernel61_Valid_Out, channel40_Kernel61_Valid_Out, channel41_Kernel61_Valid_Out, channel42_Kernel61_Valid_Out, channel43_Kernel61_Valid_Out, channel44_Kernel61_Valid_Out, channel45_Kernel61_Valid_Out, channel46_Kernel61_Valid_Out, channel47_Kernel61_Valid_Out, channel48_Kernel61_Valid_Out, channel49_Kernel61_Valid_Out, channel50_Kernel61_Valid_Out, channel51_Kernel61_Valid_Out, channel52_Kernel61_Valid_Out, channel53_Kernel61_Valid_Out, channel54_Kernel61_Valid_Out, channel55_Kernel61_Valid_Out, channel56_Kernel61_Valid_Out, channel57_Kernel61_Valid_Out, channel58_Kernel61_Valid_Out, channel59_Kernel61_Valid_Out, channel60_Kernel61_Valid_Out, channel61_Kernel61_Valid_Out, channel62_Kernel61_Valid_Out, channel63_Kernel61_Valid_Out, channel64_Kernel61_Valid_Out;

	assign add_kernel61=channel1_Kernel61_Valid_Out & channel2_Kernel61_Valid_Out & channel3_Kernel61_Valid_Out & channel4_Kernel61_Valid_Out & channel5_Kernel61_Valid_Out & channel6_Kernel61_Valid_Out & channel7_Kernel61_Valid_Out & channel8_Kernel61_Valid_Out & channel9_Kernel61_Valid_Out & channel10_Kernel61_Valid_Out & channel11_Kernel61_Valid_Out & channel12_Kernel61_Valid_Out & channel13_Kernel61_Valid_Out & channel14_Kernel61_Valid_Out & channel15_Kernel61_Valid_Out & channel16_Kernel61_Valid_Out & channel17_Kernel61_Valid_Out & channel18_Kernel61_Valid_Out & channel19_Kernel61_Valid_Out & channel20_Kernel61_Valid_Out & channel21_Kernel61_Valid_Out & channel22_Kernel61_Valid_Out & channel23_Kernel61_Valid_Out & channel24_Kernel61_Valid_Out & channel25_Kernel61_Valid_Out & channel26_Kernel61_Valid_Out & channel27_Kernel61_Valid_Out & channel28_Kernel61_Valid_Out & channel29_Kernel61_Valid_Out & channel30_Kernel61_Valid_Out & channel31_Kernel61_Valid_Out & channel32_Kernel61_Valid_Out & channel33_Kernel61_Valid_Out & channel34_Kernel61_Valid_Out & channel35_Kernel61_Valid_Out & channel36_Kernel61_Valid_Out & channel37_Kernel61_Valid_Out & channel38_Kernel61_Valid_Out & channel39_Kernel61_Valid_Out & channel40_Kernel61_Valid_Out & channel41_Kernel61_Valid_Out & channel42_Kernel61_Valid_Out & channel43_Kernel61_Valid_Out & channel44_Kernel61_Valid_Out & channel45_Kernel61_Valid_Out & channel46_Kernel61_Valid_Out & channel47_Kernel61_Valid_Out & channel48_Kernel61_Valid_Out & channel49_Kernel61_Valid_Out & channel50_Kernel61_Valid_Out & channel51_Kernel61_Valid_Out & channel52_Kernel61_Valid_Out & channel53_Kernel61_Valid_Out & channel54_Kernel61_Valid_Out & channel55_Kernel61_Valid_Out & channel56_Kernel61_Valid_Out & channel57_Kernel61_Valid_Out & channel58_Kernel61_Valid_Out & channel59_Kernel61_Valid_Out & channel60_Kernel61_Valid_Out & channel61_Kernel61_Valid_Out & channel62_Kernel61_Valid_Out & channel63_Kernel61_Valid_Out & channel64_Kernel61_Valid_Out;

	wire channel1_Kernel62_Valid_Out, channel2_Kernel62_Valid_Out, channel3_Kernel62_Valid_Out, channel4_Kernel62_Valid_Out, channel5_Kernel62_Valid_Out, channel6_Kernel62_Valid_Out, channel7_Kernel62_Valid_Out, channel8_Kernel62_Valid_Out, channel9_Kernel62_Valid_Out, channel10_Kernel62_Valid_Out, channel11_Kernel62_Valid_Out, channel12_Kernel62_Valid_Out, channel13_Kernel62_Valid_Out, channel14_Kernel62_Valid_Out, channel15_Kernel62_Valid_Out, channel16_Kernel62_Valid_Out, channel17_Kernel62_Valid_Out, channel18_Kernel62_Valid_Out, channel19_Kernel62_Valid_Out, channel20_Kernel62_Valid_Out, channel21_Kernel62_Valid_Out, channel22_Kernel62_Valid_Out, channel23_Kernel62_Valid_Out, channel24_Kernel62_Valid_Out, channel25_Kernel62_Valid_Out, channel26_Kernel62_Valid_Out, channel27_Kernel62_Valid_Out, channel28_Kernel62_Valid_Out, channel29_Kernel62_Valid_Out, channel30_Kernel62_Valid_Out, channel31_Kernel62_Valid_Out, channel32_Kernel62_Valid_Out, channel33_Kernel62_Valid_Out, channel34_Kernel62_Valid_Out, channel35_Kernel62_Valid_Out, channel36_Kernel62_Valid_Out, channel37_Kernel62_Valid_Out, channel38_Kernel62_Valid_Out, channel39_Kernel62_Valid_Out, channel40_Kernel62_Valid_Out, channel41_Kernel62_Valid_Out, channel42_Kernel62_Valid_Out, channel43_Kernel62_Valid_Out, channel44_Kernel62_Valid_Out, channel45_Kernel62_Valid_Out, channel46_Kernel62_Valid_Out, channel47_Kernel62_Valid_Out, channel48_Kernel62_Valid_Out, channel49_Kernel62_Valid_Out, channel50_Kernel62_Valid_Out, channel51_Kernel62_Valid_Out, channel52_Kernel62_Valid_Out, channel53_Kernel62_Valid_Out, channel54_Kernel62_Valid_Out, channel55_Kernel62_Valid_Out, channel56_Kernel62_Valid_Out, channel57_Kernel62_Valid_Out, channel58_Kernel62_Valid_Out, channel59_Kernel62_Valid_Out, channel60_Kernel62_Valid_Out, channel61_Kernel62_Valid_Out, channel62_Kernel62_Valid_Out, channel63_Kernel62_Valid_Out, channel64_Kernel62_Valid_Out;

	assign add_kernel62=channel1_Kernel62_Valid_Out & channel2_Kernel62_Valid_Out & channel3_Kernel62_Valid_Out & channel4_Kernel62_Valid_Out & channel5_Kernel62_Valid_Out & channel6_Kernel62_Valid_Out & channel7_Kernel62_Valid_Out & channel8_Kernel62_Valid_Out & channel9_Kernel62_Valid_Out & channel10_Kernel62_Valid_Out & channel11_Kernel62_Valid_Out & channel12_Kernel62_Valid_Out & channel13_Kernel62_Valid_Out & channel14_Kernel62_Valid_Out & channel15_Kernel62_Valid_Out & channel16_Kernel62_Valid_Out & channel17_Kernel62_Valid_Out & channel18_Kernel62_Valid_Out & channel19_Kernel62_Valid_Out & channel20_Kernel62_Valid_Out & channel21_Kernel62_Valid_Out & channel22_Kernel62_Valid_Out & channel23_Kernel62_Valid_Out & channel24_Kernel62_Valid_Out & channel25_Kernel62_Valid_Out & channel26_Kernel62_Valid_Out & channel27_Kernel62_Valid_Out & channel28_Kernel62_Valid_Out & channel29_Kernel62_Valid_Out & channel30_Kernel62_Valid_Out & channel31_Kernel62_Valid_Out & channel32_Kernel62_Valid_Out & channel33_Kernel62_Valid_Out & channel34_Kernel62_Valid_Out & channel35_Kernel62_Valid_Out & channel36_Kernel62_Valid_Out & channel37_Kernel62_Valid_Out & channel38_Kernel62_Valid_Out & channel39_Kernel62_Valid_Out & channel40_Kernel62_Valid_Out & channel41_Kernel62_Valid_Out & channel42_Kernel62_Valid_Out & channel43_Kernel62_Valid_Out & channel44_Kernel62_Valid_Out & channel45_Kernel62_Valid_Out & channel46_Kernel62_Valid_Out & channel47_Kernel62_Valid_Out & channel48_Kernel62_Valid_Out & channel49_Kernel62_Valid_Out & channel50_Kernel62_Valid_Out & channel51_Kernel62_Valid_Out & channel52_Kernel62_Valid_Out & channel53_Kernel62_Valid_Out & channel54_Kernel62_Valid_Out & channel55_Kernel62_Valid_Out & channel56_Kernel62_Valid_Out & channel57_Kernel62_Valid_Out & channel58_Kernel62_Valid_Out & channel59_Kernel62_Valid_Out & channel60_Kernel62_Valid_Out & channel61_Kernel62_Valid_Out & channel62_Kernel62_Valid_Out & channel63_Kernel62_Valid_Out & channel64_Kernel62_Valid_Out;

	wire channel1_Kernel63_Valid_Out, channel2_Kernel63_Valid_Out, channel3_Kernel63_Valid_Out, channel4_Kernel63_Valid_Out, channel5_Kernel63_Valid_Out, channel6_Kernel63_Valid_Out, channel7_Kernel63_Valid_Out, channel8_Kernel63_Valid_Out, channel9_Kernel63_Valid_Out, channel10_Kernel63_Valid_Out, channel11_Kernel63_Valid_Out, channel12_Kernel63_Valid_Out, channel13_Kernel63_Valid_Out, channel14_Kernel63_Valid_Out, channel15_Kernel63_Valid_Out, channel16_Kernel63_Valid_Out, channel17_Kernel63_Valid_Out, channel18_Kernel63_Valid_Out, channel19_Kernel63_Valid_Out, channel20_Kernel63_Valid_Out, channel21_Kernel63_Valid_Out, channel22_Kernel63_Valid_Out, channel23_Kernel63_Valid_Out, channel24_Kernel63_Valid_Out, channel25_Kernel63_Valid_Out, channel26_Kernel63_Valid_Out, channel27_Kernel63_Valid_Out, channel28_Kernel63_Valid_Out, channel29_Kernel63_Valid_Out, channel30_Kernel63_Valid_Out, channel31_Kernel63_Valid_Out, channel32_Kernel63_Valid_Out, channel33_Kernel63_Valid_Out, channel34_Kernel63_Valid_Out, channel35_Kernel63_Valid_Out, channel36_Kernel63_Valid_Out, channel37_Kernel63_Valid_Out, channel38_Kernel63_Valid_Out, channel39_Kernel63_Valid_Out, channel40_Kernel63_Valid_Out, channel41_Kernel63_Valid_Out, channel42_Kernel63_Valid_Out, channel43_Kernel63_Valid_Out, channel44_Kernel63_Valid_Out, channel45_Kernel63_Valid_Out, channel46_Kernel63_Valid_Out, channel47_Kernel63_Valid_Out, channel48_Kernel63_Valid_Out, channel49_Kernel63_Valid_Out, channel50_Kernel63_Valid_Out, channel51_Kernel63_Valid_Out, channel52_Kernel63_Valid_Out, channel53_Kernel63_Valid_Out, channel54_Kernel63_Valid_Out, channel55_Kernel63_Valid_Out, channel56_Kernel63_Valid_Out, channel57_Kernel63_Valid_Out, channel58_Kernel63_Valid_Out, channel59_Kernel63_Valid_Out, channel60_Kernel63_Valid_Out, channel61_Kernel63_Valid_Out, channel62_Kernel63_Valid_Out, channel63_Kernel63_Valid_Out, channel64_Kernel63_Valid_Out;

	assign add_kernel63=channel1_Kernel63_Valid_Out & channel2_Kernel63_Valid_Out & channel3_Kernel63_Valid_Out & channel4_Kernel63_Valid_Out & channel5_Kernel63_Valid_Out & channel6_Kernel63_Valid_Out & channel7_Kernel63_Valid_Out & channel8_Kernel63_Valid_Out & channel9_Kernel63_Valid_Out & channel10_Kernel63_Valid_Out & channel11_Kernel63_Valid_Out & channel12_Kernel63_Valid_Out & channel13_Kernel63_Valid_Out & channel14_Kernel63_Valid_Out & channel15_Kernel63_Valid_Out & channel16_Kernel63_Valid_Out & channel17_Kernel63_Valid_Out & channel18_Kernel63_Valid_Out & channel19_Kernel63_Valid_Out & channel20_Kernel63_Valid_Out & channel21_Kernel63_Valid_Out & channel22_Kernel63_Valid_Out & channel23_Kernel63_Valid_Out & channel24_Kernel63_Valid_Out & channel25_Kernel63_Valid_Out & channel26_Kernel63_Valid_Out & channel27_Kernel63_Valid_Out & channel28_Kernel63_Valid_Out & channel29_Kernel63_Valid_Out & channel30_Kernel63_Valid_Out & channel31_Kernel63_Valid_Out & channel32_Kernel63_Valid_Out & channel33_Kernel63_Valid_Out & channel34_Kernel63_Valid_Out & channel35_Kernel63_Valid_Out & channel36_Kernel63_Valid_Out & channel37_Kernel63_Valid_Out & channel38_Kernel63_Valid_Out & channel39_Kernel63_Valid_Out & channel40_Kernel63_Valid_Out & channel41_Kernel63_Valid_Out & channel42_Kernel63_Valid_Out & channel43_Kernel63_Valid_Out & channel44_Kernel63_Valid_Out & channel45_Kernel63_Valid_Out & channel46_Kernel63_Valid_Out & channel47_Kernel63_Valid_Out & channel48_Kernel63_Valid_Out & channel49_Kernel63_Valid_Out & channel50_Kernel63_Valid_Out & channel51_Kernel63_Valid_Out & channel52_Kernel63_Valid_Out & channel53_Kernel63_Valid_Out & channel54_Kernel63_Valid_Out & channel55_Kernel63_Valid_Out & channel56_Kernel63_Valid_Out & channel57_Kernel63_Valid_Out & channel58_Kernel63_Valid_Out & channel59_Kernel63_Valid_Out & channel60_Kernel63_Valid_Out & channel61_Kernel63_Valid_Out & channel62_Kernel63_Valid_Out & channel63_Kernel63_Valid_Out & channel64_Kernel63_Valid_Out;

	wire channel1_Kernel64_Valid_Out, channel2_Kernel64_Valid_Out, channel3_Kernel64_Valid_Out, channel4_Kernel64_Valid_Out, channel5_Kernel64_Valid_Out, channel6_Kernel64_Valid_Out, channel7_Kernel64_Valid_Out, channel8_Kernel64_Valid_Out, channel9_Kernel64_Valid_Out, channel10_Kernel64_Valid_Out, channel11_Kernel64_Valid_Out, channel12_Kernel64_Valid_Out, channel13_Kernel64_Valid_Out, channel14_Kernel64_Valid_Out, channel15_Kernel64_Valid_Out, channel16_Kernel64_Valid_Out, channel17_Kernel64_Valid_Out, channel18_Kernel64_Valid_Out, channel19_Kernel64_Valid_Out, channel20_Kernel64_Valid_Out, channel21_Kernel64_Valid_Out, channel22_Kernel64_Valid_Out, channel23_Kernel64_Valid_Out, channel24_Kernel64_Valid_Out, channel25_Kernel64_Valid_Out, channel26_Kernel64_Valid_Out, channel27_Kernel64_Valid_Out, channel28_Kernel64_Valid_Out, channel29_Kernel64_Valid_Out, channel30_Kernel64_Valid_Out, channel31_Kernel64_Valid_Out, channel32_Kernel64_Valid_Out, channel33_Kernel64_Valid_Out, channel34_Kernel64_Valid_Out, channel35_Kernel64_Valid_Out, channel36_Kernel64_Valid_Out, channel37_Kernel64_Valid_Out, channel38_Kernel64_Valid_Out, channel39_Kernel64_Valid_Out, channel40_Kernel64_Valid_Out, channel41_Kernel64_Valid_Out, channel42_Kernel64_Valid_Out, channel43_Kernel64_Valid_Out, channel44_Kernel64_Valid_Out, channel45_Kernel64_Valid_Out, channel46_Kernel64_Valid_Out, channel47_Kernel64_Valid_Out, channel48_Kernel64_Valid_Out, channel49_Kernel64_Valid_Out, channel50_Kernel64_Valid_Out, channel51_Kernel64_Valid_Out, channel52_Kernel64_Valid_Out, channel53_Kernel64_Valid_Out, channel54_Kernel64_Valid_Out, channel55_Kernel64_Valid_Out, channel56_Kernel64_Valid_Out, channel57_Kernel64_Valid_Out, channel58_Kernel64_Valid_Out, channel59_Kernel64_Valid_Out, channel60_Kernel64_Valid_Out, channel61_Kernel64_Valid_Out, channel62_Kernel64_Valid_Out, channel63_Kernel64_Valid_Out, channel64_Kernel64_Valid_Out;

	assign add_kernel64=channel1_Kernel64_Valid_Out & channel2_Kernel64_Valid_Out & channel3_Kernel64_Valid_Out & channel4_Kernel64_Valid_Out & channel5_Kernel64_Valid_Out & channel6_Kernel64_Valid_Out & channel7_Kernel64_Valid_Out & channel8_Kernel64_Valid_Out & channel9_Kernel64_Valid_Out & channel10_Kernel64_Valid_Out & channel11_Kernel64_Valid_Out & channel12_Kernel64_Valid_Out & channel13_Kernel64_Valid_Out & channel14_Kernel64_Valid_Out & channel15_Kernel64_Valid_Out & channel16_Kernel64_Valid_Out & channel17_Kernel64_Valid_Out & channel18_Kernel64_Valid_Out & channel19_Kernel64_Valid_Out & channel20_Kernel64_Valid_Out & channel21_Kernel64_Valid_Out & channel22_Kernel64_Valid_Out & channel23_Kernel64_Valid_Out & channel24_Kernel64_Valid_Out & channel25_Kernel64_Valid_Out & channel26_Kernel64_Valid_Out & channel27_Kernel64_Valid_Out & channel28_Kernel64_Valid_Out & channel29_Kernel64_Valid_Out & channel30_Kernel64_Valid_Out & channel31_Kernel64_Valid_Out & channel32_Kernel64_Valid_Out & channel33_Kernel64_Valid_Out & channel34_Kernel64_Valid_Out & channel35_Kernel64_Valid_Out & channel36_Kernel64_Valid_Out & channel37_Kernel64_Valid_Out & channel38_Kernel64_Valid_Out & channel39_Kernel64_Valid_Out & channel40_Kernel64_Valid_Out & channel41_Kernel64_Valid_Out & channel42_Kernel64_Valid_Out & channel43_Kernel64_Valid_Out & channel44_Kernel64_Valid_Out & channel45_Kernel64_Valid_Out & channel46_Kernel64_Valid_Out & channel47_Kernel64_Valid_Out & channel48_Kernel64_Valid_Out & channel49_Kernel64_Valid_Out & channel50_Kernel64_Valid_Out & channel51_Kernel64_Valid_Out & channel52_Kernel64_Valid_Out & channel53_Kernel64_Valid_Out & channel54_Kernel64_Valid_Out & channel55_Kernel64_Valid_Out & channel56_Kernel64_Valid_Out & channel57_Kernel64_Valid_Out & channel58_Kernel64_Valid_Out & channel59_Kernel64_Valid_Out & channel60_Kernel64_Valid_Out & channel61_Kernel64_Valid_Out & channel62_Kernel64_Valid_Out & channel63_Kernel64_Valid_Out & channel64_Kernel64_Valid_Out;


	wire [31:0] bn1_Data_Out, bn2_Data_Out, bn3_Data_Out, bn4_Data_Out, bn5_Data_Out, bn6_Data_Out, bn7_Data_Out, bn8_Data_Out, bn9_Data_Out, bn10_Data_Out, bn11_Data_Out, bn12_Data_Out, bn13_Data_Out, bn14_Data_Out, bn15_Data_Out, bn16_Data_Out, bn17_Data_Out, bn18_Data_Out, bn19_Data_Out, bn20_Data_Out, bn21_Data_Out, bn22_Data_Out, bn23_Data_Out, bn24_Data_Out, bn25_Data_Out, bn26_Data_Out, bn27_Data_Out, bn28_Data_Out, bn29_Data_Out, bn30_Data_Out, bn31_Data_Out, bn32_Data_Out, bn33_Data_Out, bn34_Data_Out, bn35_Data_Out, bn36_Data_Out, bn37_Data_Out, bn38_Data_Out, bn39_Data_Out, bn40_Data_Out, bn41_Data_Out, bn42_Data_Out, bn43_Data_Out, bn44_Data_Out, bn45_Data_Out, bn46_Data_Out, bn47_Data_Out, bn48_Data_Out, bn49_Data_Out, bn50_Data_Out, bn51_Data_Out, bn52_Data_Out, bn53_Data_Out, bn54_Data_Out, bn55_Data_Out, bn56_Data_Out, bn57_Data_Out, bn58_Data_Out, bn59_Data_Out, bn60_Data_Out, bn61_Data_Out, bn62_Data_Out, bn63_Data_Out, bn64_Data_Out;

	wire bn1_Valid_Out, bn2_Valid_Out, bn3_Valid_Out, bn4_Valid_Out, bn5_Valid_Out, bn6_Valid_Out, bn7_Valid_Out, bn8_Valid_Out, bn9_Valid_Out, bn10_Valid_Out, bn11_Valid_Out, bn12_Valid_Out, bn13_Valid_Out, bn14_Valid_Out, bn15_Valid_Out, bn16_Valid_Out, bn17_Valid_Out, bn18_Valid_Out, bn19_Valid_Out, bn20_Valid_Out, bn21_Valid_Out, bn22_Valid_Out, bn23_Valid_Out, bn24_Valid_Out, bn25_Valid_Out, bn26_Valid_Out, bn27_Valid_Out, bn28_Valid_Out, bn29_Valid_Out, bn30_Valid_Out, bn31_Valid_Out, bn32_Valid_Out, bn33_Valid_Out, bn34_Valid_Out, bn35_Valid_Out, bn36_Valid_Out, bn37_Valid_Out, bn38_Valid_Out, bn39_Valid_Out, bn40_Valid_Out, bn41_Valid_Out, bn42_Valid_Out, bn43_Valid_Out, bn44_Valid_Out, bn45_Valid_Out, bn46_Valid_Out, bn47_Valid_Out, bn48_Valid_Out, bn49_Valid_Out, bn50_Valid_Out, bn51_Valid_Out, bn52_Valid_Out, bn53_Valid_Out, bn54_Valid_Out, bn55_Valid_Out, bn56_Valid_Out, bn57_Valid_Out, bn58_Valid_Out, bn59_Valid_Out, bn60_Valid_Out, bn61_Valid_Out, bn62_Valid_Out, bn63_Valid_Out, bn64_Valid_Out;

	wire rl1_Valid_Out, rl2_Valid_Out, rl3_Valid_Out, rl4_Valid_Out, rl5_Valid_Out, rl6_Valid_Out, rl7_Valid_Out, rl8_Valid_Out, rl9_Valid_Out, rl10_Valid_Out, rl11_Valid_Out, rl12_Valid_Out, rl13_Valid_Out, rl14_Valid_Out, rl15_Valid_Out, rl16_Valid_Out, rl17_Valid_Out, rl18_Valid_Out, rl19_Valid_Out, rl20_Valid_Out, rl21_Valid_Out, rl22_Valid_Out, rl23_Valid_Out, rl24_Valid_Out, rl25_Valid_Out, rl26_Valid_Out, rl27_Valid_Out, rl28_Valid_Out, rl29_Valid_Out, rl30_Valid_Out, rl31_Valid_Out, rl32_Valid_Out, rl33_Valid_Out, rl34_Valid_Out, rl35_Valid_Out, rl36_Valid_Out, rl37_Valid_Out, rl38_Valid_Out, rl39_Valid_Out, rl40_Valid_Out, rl41_Valid_Out, rl42_Valid_Out, rl43_Valid_Out, rl44_Valid_Out, rl45_Valid_Out, rl46_Valid_Out, rl47_Valid_Out, rl48_Valid_Out, rl49_Valid_Out, rl50_Valid_Out, rl51_Valid_Out, rl52_Valid_Out, rl53_Valid_Out, rl54_Valid_Out, rl55_Valid_Out, rl56_Valid_Out, rl57_Valid_Out, rl58_Valid_Out, rl59_Valid_Out, rl60_Valid_Out, rl61_Valid_Out, rl62_Valid_Out, rl63_Valid_Out, rl64_Valid_Out;

	 assign Valid_Out = rl1_Valid_Out & rl2_Valid_Out & rl3_Valid_Out & rl4_Valid_Out & rl5_Valid_Out & rl6_Valid_Out & rl7_Valid_Out & rl8_Valid_Out & rl9_Valid_Out & rl10_Valid_Out & rl11_Valid_Out & rl12_Valid_Out & rl13_Valid_Out & rl14_Valid_Out & rl15_Valid_Out & rl16_Valid_Out & rl17_Valid_Out & rl18_Valid_Out & rl19_Valid_Out & rl20_Valid_Out & rl21_Valid_Out & rl22_Valid_Out & rl23_Valid_Out & rl24_Valid_Out & rl25_Valid_Out & rl26_Valid_Out & rl27_Valid_Out & rl28_Valid_Out & rl29_Valid_Out & rl30_Valid_Out & rl31_Valid_Out & rl32_Valid_Out & rl33_Valid_Out & rl34_Valid_Out & rl35_Valid_Out & rl36_Valid_Out & rl37_Valid_Out & rl38_Valid_Out & rl39_Valid_Out & rl40_Valid_Out & rl41_Valid_Out & rl42_Valid_Out & rl43_Valid_Out & rl44_Valid_Out & rl45_Valid_Out & rl46_Valid_Out & rl47_Valid_Out & rl48_Valid_Out & rl49_Valid_Out & rl50_Valid_Out & rl51_Valid_Out & rl52_Valid_Out & rl53_Valid_Out & rl54_Valid_Out & rl55_Valid_Out & rl56_Valid_Out & rl57_Valid_Out & rl58_Valid_Out & rl59_Valid_Out & rl60_Valid_Out & rl61_Valid_Out & rl62_Valid_Out & rl63_Valid_Out & rl64_Valid_Out;
//////////KERNEL1//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111101010001100001110001110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111110011001110110111111100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110000110111011000011000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111101111001010011001100011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111110101100000011000100111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111100100100011100101100110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111110100101111001111111100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111110111000101100110111111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111110011000000111011100001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111101100001101100000001111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111110011010110001001001101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111111000011001100111110100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111111000010000010100001000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111110011010101010101101001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110001001011100011001001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111111001111000011010011101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110101110000100111011010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110111110100100011000111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110010100111100011010010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110101111000001111111001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111111000001011101001011001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111110110110010001100001101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111110000000000100101010111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111110010100011010100111010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111110100000101011100010100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111111001000100001000110011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111111000100010110111101111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111110111000110101000100110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111110110101000110100010011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110000101100000001100111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111101100110000010010011001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111110110100101011110101010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b00111101100100011010101011101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111101101000000110011100111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111110100011100110110111000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111110100101000010001100101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b10111110010101100100110011000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111100111100001001111000100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b00111110011000111011111010101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b00111110101000011011100110010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111110010110011010100110000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111110000010110011011110011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111100010010011011011101100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b00111101100111110001011001001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111101110010100101000000000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b10111110110111001100001101100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b10111110100011101010101101011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b00111101011011011110011101010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b00111101110011010110100100111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111110111010000100011110001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b10111101110010101100111001100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111101110001000111100001000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b00111111011110010000001100011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111111001001101110011011000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111110101010111100000001101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111111100110101111111110011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b10111110110011100000100111111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b10111110001001010100111011111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b10111110110100110111101111010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b00111110011000111011010011101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b10111101110101001101100100000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b10111110101000011101001000111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b10111110011100011100001000001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111101100110101011111111110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel1_Valid_Out)
	);
	Adder_64input add_k1(
		.Data1(Data_Out_Kernel1[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel1[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel1[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel1[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel1[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel1[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel1[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel1[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel1[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel1[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel1[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel1[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel1[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel1[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel1[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel1[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel1[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel1[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel1[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel1[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel1[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel1[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel1[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel1[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel1[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel1[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel1[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel1[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel1[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel1[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel1[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel1[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel1[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel1[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel1[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel1[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel1[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel1[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel1[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel1[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel1[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel1[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel1[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel1[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel1[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel1[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel1[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel1[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel1[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel1[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel1[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel1[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel1[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel1[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel1[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel1[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel1[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel1[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel1[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel1[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel1[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel1[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel1[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel1[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel1),
		.Data_Out(add_k1_Data_Out),
		.Valid_Out(add_kernel1_Valid_Out)
	);
	Batch_Norm bn_kernel1(
		.Data_A(32'b00111110110101000111000000001111),
		.Data_B(32'b00111111011101011100010110000111),
		.Data_In(add_k1_Data_Out),
		.Valid_In(add_kernel1_Valid_Out),
		.Data_Out(bn1_Data_Out),
		.Valid_Out(bn1_Valid_Out)
	);
	Relu_Core rl_kernel1(
		.Data_In(bn1_Data_Out),
		.Valid_In(bn1_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT-1:0]),
		.Valid_Out(rl1_Valid_Out)
	);
//////////KERNEL2//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111110000011001110000010001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110111111110101101010101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110101010111000011010010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111111100001000100011000001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111101100111011101111101111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111101101101110010100010101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111110101110101100101000110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111011001101000000001111111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111110110001100101010100011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111110011100010011011001101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110011000111000011000000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111110100101001000011000010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110110101110001110011000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111110110101100101000001101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110101010000100010101001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111110110010100000111010000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110000000011001111000101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111011111001001101111010110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110100101110001111100101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111011010111000011110011100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110110101101011101110101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111101110111001101110111100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111110101100000000001011010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111111010101001111001110110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111111000010111101011001011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111111010011010110011101011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110101011100101100010001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111101110010010010110100101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111111000011111110010110110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111101100111111111000010000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111110111010000011110111011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111101110111010011011111110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111101111011111100100101111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111110101101010010010100011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111110000110110000110000101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b10111100111000011110101100010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111101101011001101111111111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b00111110010001101011000111101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111101111110001111001000101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b00111110111011110011010011000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111110100111001111011001110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111111000011110111111001001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111111001001010111101101001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b00111110100101101010101110001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b00111110011110111110000001110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b10111101111101110001111110100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b10111110001011010110011000000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111100110101011011100000111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111101101110101100100111000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b00111110000011011010000001100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111111000010101110010101010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111110110110110110110010001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111110011111011011110011011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b00111110111011111101100001101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111110100100000001000001000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b00111110101110000010000001010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b10111110111000101001011011010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111111000100000100001001111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b10111110110100100101111011001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b00111110000111011100000001000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111101001111001011110101111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111110100001100011010111011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b10111100011111001100010101101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b10111110110000010000010011110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel2_Valid_Out)
	);
	Adder_64input add_k2(
		.Data1(Data_Out_Kernel2[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel2[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel2[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel2[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel2[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel2[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel2[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel2[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel2[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel2[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel2[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel2[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel2[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel2[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel2[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel2[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel2[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel2[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel2[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel2[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel2[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel2[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel2[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel2[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel2[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel2[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel2[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel2[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel2[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel2[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel2[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel2[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel2[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel2[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel2[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel2[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel2[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel2[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel2[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel2[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel2[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel2[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel2[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel2[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel2[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel2[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel2[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel2[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel2[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel2[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel2[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel2[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel2[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel2[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel2[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel2[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel2[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel2[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel2[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel2[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel2[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel2[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel2[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel2[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel2),
		.Data_Out(add_k2_Data_Out),
		.Valid_Out(add_kernel2_Valid_Out)
	);
	Batch_Norm bn_kernel2(
		.Data_A(32'b00111110111000011011011011110100),
		.Data_B(32'b00111111010010111101011100110010),
		.Data_In(add_k2_Data_Out),
		.Valid_In(add_kernel2_Valid_Out),
		.Data_Out(bn2_Data_Out),
		.Valid_Out(bn2_Valid_Out)
	);
	Relu_Core rl_kernel2(
		.Data_In(bn2_Data_Out),
		.Valid_In(bn2_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Valid_Out(rl2_Valid_Out)
	);
//////////KERNEL3//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111111000111101001000110011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110111000011110111111000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110001111101000100011010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110001101111000101000100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111101110111100001110001001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111110011000000100110011011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111111000010010111110000000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111101001101011110110100010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110000110110111011111110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111110101100010010010001101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111101010011101110011011001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111111010000010111001110001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110001010000010011011011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111110100000000010111110000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110001001110000001011001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111110100001010111100001101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110010000011000111001101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111101100110101001011111000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111101001100011101111010100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110001010000001001001001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110010110101110110100111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111110010011010001001110110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111101100011010100010110111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111110111111010111110011100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111110101100111100000011010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110101110010000110011100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110110001011000000010100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111110011110000011101111000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111111010011110011001100000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111100100100011111000110110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111110110101101000111010110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111111001000000100110011010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111100011110010011001001011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111110111000001110100010111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111110111100101101101000010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111110001000000010001111000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b10111100110011100110100100100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111110100001011111100010111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b00111110000110011101001100010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111111001101011001110000111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111111011000100000100110101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111110001110100111100101100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b00111100001100100010000101011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111101111011011001000101110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b00111110100011110101010010011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111111000111111100010011000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b10111110101010001000010110010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111110110111100010010110001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111101000111011000011111010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111111000010001001010111101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111101000101101011000101010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111110000101110111010111000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b00111110110101001100001010110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b00111110010010000001110010000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111111000110001111100000111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111110100001001111111110000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111101101001100000011011111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b10111110101011000100111111010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b10111110111101011111000001000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111110101111101000110101001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111110101000001011101011110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b10111110110101010100100111011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b10111111011110100101110111111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b10111110111100101010000010100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel3_Valid_Out)
	);
	Adder_64input add_k3(
		.Data1(Data_Out_Kernel3[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel3[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel3[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel3[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel3[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel3[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel3[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel3[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel3[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel3[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel3[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel3[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel3[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel3[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel3[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel3[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel3[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel3[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel3[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel3[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel3[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel3[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel3[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel3[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel3[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel3[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel3[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel3[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel3[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel3[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel3[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel3[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel3[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel3[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel3[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel3[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel3[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel3[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel3[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel3[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel3[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel3[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel3[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel3[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel3[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel3[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel3[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel3[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel3[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel3[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel3[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel3[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel3[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel3[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel3[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel3[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel3[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel3[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel3[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel3[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel3[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel3[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel3[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel3[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel3),
		.Data_Out(add_k3_Data_Out),
		.Valid_Out(add_kernel3_Valid_Out)
	);
	Batch_Norm bn_kernel3(
		.Data_A(32'b00111110110111110111100111110001),
		.Data_B(32'b00111111010111001001111101001001),
		.Data_In(add_k3_Data_Out),
		.Valid_In(add_kernel3_Valid_Out),
		.Data_Out(bn3_Data_Out),
		.Valid_Out(bn3_Valid_Out)
	);
	Relu_Core rl_kernel3(
		.Data_In(bn3_Data_Out),
		.Valid_In(bn3_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(rl3_Valid_Out)
	);
//////////KERNEL4//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111101010110010001011000011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111101001001000100101110110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110101011100100011011100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110101011101001010101111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111110000011001011010100111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111110000100110001110111100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111111000100010110001111100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111110111101000001101000100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111111001010110101000011011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111110101001010101000110100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111111000011110111010010010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111110111000100010001001001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111111000010000110111110100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111110001101011111110000010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111111000110010111011110100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111101100011111110000101001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111110111101111000000101011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111110010000111000000001110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111111001010011111100101110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110010101111100000111101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110100011000000101000101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111110101111110011110110000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111110101111111110111000100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111110000110101110000000100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111110100110111001010100001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111110111001101001111000000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111110011110101001010000100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111110000100100101011000011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111101100011101001000001101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111101100110001101101111011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111111001110101111100000110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110100111110010000001101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b00111101111100110100000010111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b00111111000100011100100101100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111110111010110001010010011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b10111110111101010011001001111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b10111110101001110111011111101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b00111110100100011011111000000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b00111101110001001100101010010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b00111101100100001001101000011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b10111101100100111100101011100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111101100000000011000110011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b00111110011100000010000011011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b00111110001000001101100100001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111110100111100101001011000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111110111001011110100011100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111101010110010111100011000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111110101000111000000000011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b00111110000110111111010001000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111110110111110101110011110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111111001010111010001011000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111110010001101100101001001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b00111101101111001000011100010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111110101111001111001111001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111110001111001101010000000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111110101010000100110110100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b10111111011001001000010100011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b10111110011101111000010110110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b10111110011111100101000110111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b00111110110111000101001110001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111110001101010001011100101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111110110000001011100110101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111110111010101101110000010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b10111100010110001010100100100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel4_Valid_Out)
	);
	Adder_64input add_k4(
		.Data1(Data_Out_Kernel4[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel4[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel4[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel4[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel4[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel4[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel4[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel4[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel4[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel4[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel4[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel4[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel4[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel4[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel4[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel4[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel4[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel4[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel4[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel4[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel4[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel4[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel4[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel4[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel4[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel4[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel4[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel4[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel4[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel4[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel4[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel4[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel4[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel4[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel4[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel4[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel4[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel4[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel4[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel4[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel4[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel4[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel4[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel4[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel4[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel4[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel4[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel4[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel4[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel4[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel4[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel4[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel4[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel4[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel4[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel4[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel4[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel4[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel4[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel4[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel4[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel4[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel4[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel4[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel4),
		.Data_Out(add_k4_Data_Out),
		.Valid_Out(add_kernel4_Valid_Out)
	);
	Batch_Norm bn_kernel4(
		.Data_A(32'b00111110110111010011110001001111),
		.Data_B(32'b00111101111100110001110001110100),
		.Data_In(add_k4_Data_Out),
		.Valid_In(add_kernel4_Valid_Out),
		.Data_Out(bn4_Data_Out),
		.Valid_Out(bn4_Valid_Out)
	);
	Relu_Core rl_kernel4(
		.Data_In(bn4_Data_Out),
		.Valid_In(bn4_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(rl4_Valid_Out)
	);
//////////KERNEL5//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111111100111110111111010101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111111001100111001111010100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110011010011011001110010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111101111101001011000101000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111110111110000100011000011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111110100111100110011100000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111110110000011010101010110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111100000010010111100111011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111111001011100001011101111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110010100011011111111011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110101011110011100110001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111111001101111011100001011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111101101111101111011111001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111101001110000010000001011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110101110011010001111001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111110000010110100000100111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110011111000010000100000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111110010011111111110100100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110010010011001000100101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111100010010110000110101001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111101011111100111010100001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111110001110011100111111011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111111001000001101100001001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111111010001011110100010101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111110101000011100110010101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110001101000010010010010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111110100010100100010011101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110000101101011110111110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111110011100011111101110011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110000110101010011100101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111110011001000011110001011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111111000011111111001100111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111101001101101100110001001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111110010111000000011101100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111110001001001111010110001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b10111110010101101001000010001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b10111110111010100010000111011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b00111111001000010101000010000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b00111011001000001011111101111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b00111110101100011110000110111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111111000000000111000011100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111100100110110101110111111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111101001110000110101101011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b00111101100000011010000100000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b00111110101011010001011101000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111110000011111110101111011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b10111011101100000010110100110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111101011111110100010110001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111110010011011110000010011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b00111100100011010001101001110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b10111111001001010001111011000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111100011001100111011111010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111100000101001010011110110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b00111101100010010010001100011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b10111110100101001010101000011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b00111110001011111111011111101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b10111110111110011011111101100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111110001111101110010000101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b10111111001101110101110011011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b00111110000011001101001100100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b10111111010100010101010110000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b10111111000001010001100110100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111110010011010001010000010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111110011000110101100110000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel5_Valid_Out)
	);
	Adder_64input add_k5(
		.Data1(Data_Out_Kernel5[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel5[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel5[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel5[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel5[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel5[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel5[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel5[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel5[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel5[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel5[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel5[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel5[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel5[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel5[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel5[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel5[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel5[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel5[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel5[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel5[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel5[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel5[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel5[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel5[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel5[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel5[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel5[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel5[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel5[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel5[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel5[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel5[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel5[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel5[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel5[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel5[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel5[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel5[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel5[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel5[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel5[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel5[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel5[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel5[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel5[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel5[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel5[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel5[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel5[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel5[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel5[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel5[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel5[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel5[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel5[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel5[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel5[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel5[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel5[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel5[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel5[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel5[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel5[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel5),
		.Data_Out(add_k5_Data_Out),
		.Valid_Out(add_kernel5_Valid_Out)
	);
	Batch_Norm bn_kernel5(
		.Data_A(32'b00111110111001011100101001110000),
		.Data_B(32'b00111111001101011101111011110001),
		.Data_In(add_k5_Data_Out),
		.Valid_In(add_kernel5_Valid_Out),
		.Data_Out(bn5_Data_Out),
		.Valid_Out(bn5_Valid_Out)
	);
	Relu_Core rl_kernel5(
		.Data_In(bn5_Data_Out),
		.Valid_In(bn5_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(rl5_Valid_Out)
	);
//////////KERNEL6//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111111010000110011001001011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111101100111001011111110001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110010100010111010101111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111101110010011110010110111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111111001001110010100111111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111111010011110101101101100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111110011100111010111111100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111111001010101000101011110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110101011011001101001100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111110100101111110100010000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111110101000100010111010011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110001000110010001011100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110101010001001101011001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111110110101111100011010011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110010000110110100100000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111011111110001101111100100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110010101000101100001011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110110111001000000011110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110111001010100000100010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110010001000100100001110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111100100110110110001011011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111100010011000010101000011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110010010101110100000101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111111000110100100100011011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111110011110011110001101111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111111000101110001000101001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111110011101110000000001010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110101011011101000010110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111111000000001011100010000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111100010001110010010111001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111110110011100010101101111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111101011011001111101111101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111110101101101011110011111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b00111101110011011010011111000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111110011010000111011111110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b10111110110110111100001010001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b10111100010010000001101101111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b00111110100111010100101100101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b00111110100001000111010101100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111110010000101101000001010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111110101101111100110100110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111110010000010111111101100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111110101011101110111111111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111110100011101000100110111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b00111110000101101111101010000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111110101010101110010001100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111110110111101010011111000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b00111110111100001000011100011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b00111111000001000000101001101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111110001011100110010010001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b10111110100111000001110011111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111110010001000110101101110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111101110010011110110101100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111110001000100010001100011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b10111110010100110110100000000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111101110010000001101100010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111110010110100000000100010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111111010000100101000111001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b10111111001111101110110000001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111110010111110000101001001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111101110111101111010111100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111110000101001110010011010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111110110101001111001000101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111110110000100000001001001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel6_Valid_Out)
	);
	Adder_64input add_k6(
		.Data1(Data_Out_Kernel6[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel6[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel6[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel6[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel6[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel6[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel6[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel6[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel6[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel6[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel6[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel6[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel6[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel6[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel6[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel6[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel6[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel6[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel6[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel6[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel6[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel6[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel6[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel6[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel6[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel6[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel6[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel6[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel6[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel6[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel6[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel6[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel6[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel6[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel6[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel6[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel6[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel6[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel6[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel6[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel6[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel6[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel6[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel6[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel6[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel6[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel6[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel6[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel6[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel6[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel6[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel6[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel6[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel6[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel6[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel6[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel6[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel6[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel6[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel6[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel6[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel6[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel6[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel6[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel6),
		.Data_Out(add_k6_Data_Out),
		.Valid_Out(add_kernel6_Valid_Out)
	);
	Batch_Norm bn_kernel6(
		.Data_A(32'b00111111000000001011011010101011),
		.Data_B(32'b10111101010000100010010111010100),
		.Data_In(add_k6_Data_Out),
		.Valid_In(add_kernel6_Valid_Out),
		.Data_Out(bn6_Data_Out),
		.Valid_Out(bn6_Valid_Out)
	);
	Relu_Core rl_kernel6(
		.Data_In(bn6_Data_Out),
		.Valid_In(bn6_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(rl6_Valid_Out)
	);
//////////KERNEL7//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110001000101001110010110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110011001000101011010001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110010111000101000001010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111111000011100111110100000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111111000100110010101111111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111101011010111011110110111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111111000011001000111000101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111110101111001100101110110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111110110001000110111101111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110010101011001111001110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110100110001100101010100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110011111100111010001000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111110111101000000100111101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111101100101000111111010010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110110110100001001001101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111101100101100100011000000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110010000000110000111101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111011110111111111100101101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110110110010100111000101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111011001000101011000111101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110100001011111001100010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111010111110001110111111001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111110001000100100101010101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111111000100001100010111110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111110010111101000000001111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111111011011011101111111110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111111000100101111011011000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110100111101010101000011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111101000010110011100101000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111110100010100011110100110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111110011110100010101010110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110010100010010100011010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111110011010110100110101101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111110000010101110001001011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111110011011010100100010110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111110101011010101011000111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111110010001101100011001100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b00111100110110011001100110101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111110110111010100001001000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b00111110001101010111110000001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111110110101100001110011011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111111001011011010111010000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111110111111110011001111011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b00111110011101100000101011001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b00111110101110011010110011101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111110010101100110001011100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111111010001010001111010101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111100010010001110010111010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111110111110111111011010111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111110011000110001000101100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111111000100111011001000011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b10111110010111111001110001110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111110101001110000001111110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111110011111001100100000011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111110111010100011110001001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b00111111010101010011110000001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111101000101011000010000000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111011010010000100011110100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111110010001101101001110000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111110111010101111101011110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b10111100100010010010110011000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b10111101010110111010101111111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111110010001110100101111111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111101101101111110010100010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel7_Valid_Out)
	);
	Adder_64input add_k7(
		.Data1(Data_Out_Kernel7[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel7[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel7[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel7[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel7[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel7[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel7[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel7[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel7[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel7[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel7[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel7[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel7[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel7[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel7[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel7[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel7[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel7[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel7[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel7[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel7[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel7[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel7[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel7[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel7[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel7[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel7[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel7[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel7[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel7[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel7[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel7[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel7[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel7[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel7[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel7[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel7[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel7[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel7[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel7[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel7[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel7[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel7[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel7[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel7[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel7[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel7[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel7[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel7[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel7[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel7[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel7[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel7[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel7[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel7[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel7[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel7[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel7[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel7[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel7[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel7[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel7[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel7[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel7[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel7),
		.Data_Out(add_k7_Data_Out),
		.Valid_Out(add_kernel7_Valid_Out)
	);
	Batch_Norm bn_kernel7(
		.Data_A(32'b00111110111001000101100101011100),
		.Data_B(32'b00111110111101100010100110100011),
		.Data_In(add_k7_Data_Out),
		.Valid_In(add_kernel7_Valid_Out),
		.Data_Out(bn7_Data_Out),
		.Valid_Out(bn7_Valid_Out)
	);
	Relu_Core rl_kernel7(
		.Data_In(bn7_Data_Out),
		.Valid_In(bn7_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(rl7_Valid_Out)
	);
//////////KERNEL8//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111101110010001010010101000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111101010111101111011111000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110110111111101101111111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110110001111010001001100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111110101110000000010110010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111101011111001001110001001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111110110100010010101111011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111110000111000110110111010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111111010111110100001000011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110110101110010011101110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110100011001110010111000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111111011110000111011101100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111110100101101110110011000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111111000001100101110011011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111011100110101111110111100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111111001010111100011000011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111111000001010111001011101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111110100001100101000110111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111110110011010011100100010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111101110010010110001001000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110000110010110000101100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111110000110100111111000100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110111101000010101001001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111101010001010110110001110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111110101111110111011100101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111101100100000011011111000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110001110110110110110111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110000001010110100011110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111111000000000101100011111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111101111101001011010010011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111100110001100111000010100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111011101111011101001011111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111101001101001111000000111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111110111101000001000001110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111110001111010011010000011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111111000000010111110001001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111100101001010111011000000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111110110011011111101101000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111110100110110001001010110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b00111101101111110010110110010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111110000100100000111101100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b10111111000011110111100110010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111110011100110110010101101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111110100111111100011100000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b00111110100010010001001011001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111110001011000001111110001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b10111101111001011000111011111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111111000100110010110101100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b00111110011100111011100110001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b00111101011110000001011010101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b10111110100011011000010011110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111101010011011101010011111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b00111111001000001101100110000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111101111000011011011101111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111111000011101110100000100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b00111110000011000110100100001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b10111111001011000000000111110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b10111110001100101010100111110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111101110111110011101001110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b00111110000000101011001001000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b10111110101100000001110001111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b10111111001011100000011001100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b10111110101010100000011100101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b10111110010010110010000100001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel8_Valid_Out)
	);
	Adder_64input add_k8(
		.Data1(Data_Out_Kernel8[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel8[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel8[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel8[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel8[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel8[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel8[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel8[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel8[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel8[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel8[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel8[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel8[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel8[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel8[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel8[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel8[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel8[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel8[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel8[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel8[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel8[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel8[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel8[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel8[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel8[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel8[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel8[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel8[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel8[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel8[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel8[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel8[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel8[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel8[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel8[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel8[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel8[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel8[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel8[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel8[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel8[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel8[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel8[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel8[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel8[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel8[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel8[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel8[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel8[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel8[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel8[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel8[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel8[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel8[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel8[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel8[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel8[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel8[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel8[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel8[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel8[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel8[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel8[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel8),
		.Data_Out(add_k8_Data_Out),
		.Valid_Out(add_kernel8_Valid_Out)
	);
	Batch_Norm bn_kernel8(
		.Data_A(32'b00111110111101000000011011111001),
		.Data_B(32'b00111110111010111111100001111000),
		.Data_In(add_k8_Data_Out),
		.Valid_In(add_kernel8_Valid_Out),
		.Data_Out(bn8_Data_Out),
		.Valid_Out(bn8_Valid_Out)
	);
	Relu_Core rl_kernel8(
		.Data_In(bn8_Data_Out),
		.Valid_In(bn8_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(rl8_Valid_Out)
	);
//////////KERNEL9//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111101110010110010111011101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111100110001001101000100110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110000110111000110101011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110010101001001001111100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111110010111010001010000000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111111001010001010011110101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111111001101110110001100111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111110011110101110011100111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110010000001110011011010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111111000000011010100100110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111110110000110110100110100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110111001010100100111111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111111000111010100000101010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111101110111000001101110000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111101001000000010100101000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111111010000001110001111000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110010001011110010010000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111110000001000001011110000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111110110010001100100010000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110110011000101100100110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111101110001001100110001000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111111000101010010000000111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111110100111011011001001010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111110011111000000001111111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111110100000100000011011001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111101010110110010000010001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111101100101010101111001000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110111011100101110010111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111111001000111111111101110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111111011010101001101101101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111110001101100011101100100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111101010101001011110101101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b00111101110011110100011001000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111111001000010110010111001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111110010111111000110001111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b10111101011110101001000111000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111110011010101100111110111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b00111110000011000001111111000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111111000000010110110000001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111110111001011011111110011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b10111111001011101011001011000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b10111110101010011111001111111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111101100011010011111100000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111100110100110010001001011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111110000000011011110100101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b10111110000101001100001110001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111110010101100010100010011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111101011010010100110011110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b00111110101100111000000111111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111111000101101110000000001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b10111111000010001000100100101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111110101100000000000001110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b00111110101000011101101101011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111100101100100010111010010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111110101101100010011001101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111101010111101001001101101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111110101000101000110000110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b10111110001110010111110000101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111110100001001000101010000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b00111110001101101010111001001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111110001111010100010000110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b10111101101000001000001100111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111101001111111011110000000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111110100111011110000000001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel9_Valid_Out)
	);
	Adder_64input add_k9(
		.Data1(Data_Out_Kernel9[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel9[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel9[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel9[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel9[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel9[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel9[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel9[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel9[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel9[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel9[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel9[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel9[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel9[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel9[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel9[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel9[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel9[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel9[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel9[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel9[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel9[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel9[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel9[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel9[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel9[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel9[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel9[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel9[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel9[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel9[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel9[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel9[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel9[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel9[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel9[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel9[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel9[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel9[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel9[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel9[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel9[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel9[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel9[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel9[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel9[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel9[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel9[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel9[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel9[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel9[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel9[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel9[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel9[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel9[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel9[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel9[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel9[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel9[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel9[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel9[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel9[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel9[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel9[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel9),
		.Data_Out(add_k9_Data_Out),
		.Valid_Out(add_kernel9_Valid_Out)
	);
	Batch_Norm bn_kernel9(
		.Data_A(32'b00111110111010001001010000110010),
		.Data_B(32'b10111110011000001011111000111010),
		.Data_In(add_k9_Data_Out),
		.Valid_In(add_kernel9_Valid_Out),
		.Data_Out(bn9_Data_Out),
		.Valid_Out(bn9_Valid_Out)
	);
	Relu_Core rl_kernel9(
		.Data_In(bn9_Data_Out),
		.Valid_In(bn9_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(rl9_Valid_Out)
	);
//////////KERNEL10//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110000001011001000011101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111101000100010011001100111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110100000011001111010100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110101111001110101000011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111100111011111011100000010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110111000000111001000100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111110000010110110000000001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111110010000001110000101011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110111100111010000100100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110100000000001110101000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111111001101111110111011101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111110010001100111100101010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110110010001000100000001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111101000010001100110111010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110100100101010010000000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111110010101011010100100110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111111001111101100011111110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110011110110111011001100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111110000011100000110010000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110100100000001100100111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111111000011110000111101110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111110000001001110011000000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110100100010101111110101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111110100000011111101101011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111110011010011011101000100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111101010001010101101111011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111110110000000001101100111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110010110010001010101101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111100101000010011110110010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110100011011110100010111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111110010000011101000110001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111111010011110010100011001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111110010001001011111110101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111111001011000011111000001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111110101001010011100111101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111110110111110010111111010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b10111100111000010011111101111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111100101011000110100000000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b00111110100001011101101011111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111110000001000111011000011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111110101001100101000001110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b10111110111000100100001011111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b00111110111110000110101101011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111110101000010101000110000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b00111110101111001000001101000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111110111001100001000000011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b10111110111011111011001000010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111111010000000000010100010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b00111110011101100011110010101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111101100101000011101101010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b10111110000111100011000001010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b10111110000110011101110111011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b00111110101101111001010011101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111110100010001011001010100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111110101010010101011110111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b00111101100111000111100011011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111110110011001000000011111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b10111111001001000110010100111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111111000110110110101100001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111110001100100100011011110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b10111100100001101110001000111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b10111110001000001101100110101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b10111101110110101100110110011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111101100010101100011101011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel10_Valid_Out)
	);
	Adder_64input add_k10(
		.Data1(Data_Out_Kernel10[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel10[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel10[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel10[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel10[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel10[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel10[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel10[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel10[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel10[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel10[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel10[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel10[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel10[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel10[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel10[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel10[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel10[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel10[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel10[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel10[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel10[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel10[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel10[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel10[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel10[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel10[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel10[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel10[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel10[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel10[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel10[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel10[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel10[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel10[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel10[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel10[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel10[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel10[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel10[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel10[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel10[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel10[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel10[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel10[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel10[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel10[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel10[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel10[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel10[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel10[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel10[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel10[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel10[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel10[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel10[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel10[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel10[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel10[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel10[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel10[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel10[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel10[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel10[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel10),
		.Data_Out(add_k10_Data_Out),
		.Valid_Out(add_kernel10_Valid_Out)
	);
	Batch_Norm bn_kernel10(
		.Data_A(32'b00111111000000011100011000111011),
		.Data_B(32'b10111110111110110000110110110101),
		.Data_In(add_k10_Data_Out),
		.Valid_In(add_kernel10_Valid_Out),
		.Data_Out(bn10_Data_Out),
		.Valid_Out(bn10_Valid_Out)
	);
	Relu_Core rl_kernel10(
		.Data_In(bn10_Data_Out),
		.Valid_In(bn10_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(rl10_Valid_Out)
	);
//////////KERNEL11//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111101101011011000001010001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110101111101010000011110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110011001001001100101111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110010110000001010011100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111110110001010010101111001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111101110000001110111100001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111100110111101100111010011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111101011110101100101100110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110001101111001011100101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110110011100000110001001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111101000010010011000001011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111111000001100010011010111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111111011000111010001110111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111101111111111011001110011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110101000101111111100110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111110010000101110110101011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110110101100000011011011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111101110100000010011100111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111101111011001101011011101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110100100010010000110111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111101111101111000010101100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111101101111101111000100100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111111000000110110100001011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111111011001110110000000000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111101011010010010110011001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111110010100001000010111001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111111000111111110010010110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111110001011110100100111011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111100111001110000010110110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111110101101010111011010111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111111000001011100001011100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111110101001101010100110110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111110010011110001011011010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111101011111011010111010010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111110000110100001001101111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111101010101100011100011000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111110111000100100111101111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111110001000101100110111111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b00111101011101111111000010101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b00111101111010110000110011111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b10111110010001110101010011011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b10111110101000111001101110101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b00111111000001000110100101101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b00111111001000111000000010011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111110101010000111101011010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111111100101001000000010101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b10111110101010100000011001010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111110100001010111111111001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111110000110001110010111111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111100011001011010000101100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111101010111011000111111000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b10111110111100001011000001001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b00111110111111101001111101001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111110110011110000101000010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111110011011001000001001111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b00111110010100100011100111010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111101111001111010111101101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b10111110010101010101010011101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111110011001011011100001100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111111001011010001001000001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111110100011000011101101110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b10111110010000011101000110111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b10111110110001101000010010111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b10111111000000110111100100111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel11_Valid_Out)
	);
	Adder_64input add_k11(
		.Data1(Data_Out_Kernel11[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel11[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel11[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel11[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel11[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel11[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel11[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel11[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel11[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel11[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel11[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel11[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel11[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel11[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel11[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel11[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel11[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel11[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel11[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel11[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel11[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel11[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel11[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel11[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel11[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel11[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel11[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel11[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel11[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel11[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel11[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel11[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel11[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel11[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel11[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel11[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel11[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel11[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel11[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel11[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel11[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel11[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel11[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel11[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel11[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel11[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel11[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel11[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel11[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel11[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel11[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel11[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel11[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel11[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel11[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel11[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel11[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel11[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel11[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel11[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel11[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel11[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel11[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel11[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel11),
		.Data_Out(add_k11_Data_Out),
		.Valid_Out(add_kernel11_Valid_Out)
	);
	Batch_Norm bn_kernel11(
		.Data_A(32'b00111110111111000000011100110101),
		.Data_B(32'b00111111000110010010011111011000),
		.Data_In(add_k11_Data_Out),
		.Valid_In(add_kernel11_Valid_Out),
		.Data_Out(bn11_Data_Out),
		.Valid_Out(bn11_Valid_Out)
	);
	Relu_Core rl_kernel11(
		.Data_In(bn11_Data_Out),
		.Valid_In(bn11_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(rl11_Valid_Out)
	);
//////////KERNEL12//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111110101010100000101001111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111110100000011011100001111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110010010101100101100110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110100001001111101011100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111111001011111111100110001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111110101001001110101100011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111110011000100110100001001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111101011011001010011110011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111011111110000111000100110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110101111110010111011001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111111010101000111000100111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111110001000011111111000101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111110110011011000010111100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111110110100100100011100110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110110000111110111110110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111100000000001011111101001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111101100100101111101111111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111101011001000010010001011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111111000011010011111010101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111101111000110111110100010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110100111011011011111101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111111010100010000001011100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111111100011000101010111011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111111000001110110000110100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111110111011100100100100010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111110110101001101111101101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111111000111100010111111111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111101100011111000001101101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111111001000111110000101111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111111001100011100100000100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111110011110100010011110101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110101000010111110010111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b00111110000011110010001110110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111101110001001101111001001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111110100101101000001100101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111110100100011100110100011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b10111101110011101101110000001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111101010110011010111000101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111110011000011000000000110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111111000011000000100000110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111110100001111100010001100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111110110110110011110001110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b00111111001100101111101001010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111111000101101110101101001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111110101011111001110110011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111101100111111111011110000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111110001011010110101100110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b00111100011110110001111100000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b00111110100111111011100110010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b00111110110010000100100001001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111110011011011101111100110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b10111100111000010110011110001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b00111101111111011101000101010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b00111110100111110101000110101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111110100100110110011011100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b00111101100000101110001110101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b10111111010010000101010000001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111101011101111011001010101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111110011001100011110001110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111101100011100110110110101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b10111110101010100100001100010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b10111110010110111011010100001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b10111010110110011010001111101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b10111110010111010101010111001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel12_Valid_Out)
	);
	Adder_64input add_k12(
		.Data1(Data_Out_Kernel12[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel12[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel12[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel12[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel12[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel12[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel12[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel12[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel12[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel12[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel12[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel12[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel12[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel12[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel12[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel12[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel12[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel12[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel12[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel12[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel12[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel12[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel12[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel12[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel12[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel12[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel12[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel12[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel12[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel12[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel12[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel12[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel12[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel12[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel12[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel12[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel12[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel12[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel12[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel12[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel12[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel12[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel12[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel12[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel12[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel12[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel12[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel12[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel12[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel12[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel12[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel12[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel12[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel12[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel12[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel12[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel12[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel12[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel12[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel12[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel12[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel12[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel12[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel12[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel12),
		.Data_Out(add_k12_Data_Out),
		.Valid_Out(add_kernel12_Valid_Out)
	);
	Batch_Norm bn_kernel12(
		.Data_A(32'b00111110111010110011001000111100),
		.Data_B(32'b00111110110101101001010110001110),
		.Data_In(add_k12_Data_Out),
		.Valid_In(add_kernel12_Valid_Out),
		.Data_Out(bn12_Data_Out),
		.Valid_Out(bn12_Valid_Out)
	);
	Relu_Core rl_kernel12(
		.Data_In(bn12_Data_Out),
		.Valid_In(bn12_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(rl12_Valid_Out)
	);
//////////KERNEL13//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111111001011011010111100111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111110001000011101000111111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111101001010000010000010001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111111011001001001000100100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111110110000110110001011011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110001001101101100000010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111110100001011110111100110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111111000010000000001110111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111110100100000100000111101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111110100001010111101100101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110000110101111000000001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111101101011101110101101101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111110100011010101000110011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111110000010000101010100111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110111000011111110011010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111111000010010000001100000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110100101011001111111010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111111010001110110111001110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111101101110111001011000100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111111000001011110111101001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111101101101100111001000110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111111010111000100110001101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110000110000011111011010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111110101001010011111001000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111111000010101010011011110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111101000010101001001100010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111101101111101111100111111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110101001010111010110110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111110111010011111100101000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111101111110001110000110100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111110100101011011100100011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110000101010011111111110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b00111110110100100011100110110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b00111110000001110101111001111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111110001001001010010001101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b10111101110010011101001010000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111110000001010101110010111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111111100100100000010001110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b00111110100101111101100011100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111011101101110000111010000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111110000001000001000111100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b10111100110101110111001111001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111101111100111110010110011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b00111110100101111001111001110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b00111101010100000110111100111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111110101100110010110001011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b10111111000100011100000100111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111110100000110010111001111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b00111110001111111101010100011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b00111110111001001110001101110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b10111111000011111001010110010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111110000111101110000110100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111110001001110000101101101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b00111100111110001100000111101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111101101000100101001000011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111011110111011110100001111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111110011101100100111010110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b10111110100000001011001101100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b10111110110100011110100110111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b00111110111111000111001001101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b10111100010100101110001101011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111110101101000010000000110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b10111110101110110010010011101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b10111110101111100010001001011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel13_Valid_Out)
	);
	Adder_64input add_k13(
		.Data1(Data_Out_Kernel13[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel13[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel13[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel13[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel13[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel13[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel13[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel13[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel13[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel13[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel13[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel13[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel13[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel13[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel13[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel13[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel13[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel13[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel13[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel13[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel13[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel13[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel13[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel13[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel13[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel13[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel13[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel13[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel13[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel13[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel13[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel13[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel13[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel13[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel13[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel13[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel13[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel13[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel13[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel13[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel13[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel13[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel13[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel13[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel13[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel13[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel13[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel13[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel13[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel13[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel13[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel13[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel13[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel13[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel13[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel13[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel13[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel13[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel13[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel13[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel13[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel13[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel13[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel13[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel13),
		.Data_Out(add_k13_Data_Out),
		.Valid_Out(add_kernel13_Valid_Out)
	);
	Batch_Norm bn_kernel13(
		.Data_A(32'b00111110110100111101101001011111),
		.Data_B(32'b00111111001100100001001101011110),
		.Data_In(add_k13_Data_Out),
		.Valid_In(add_kernel13_Valid_Out),
		.Data_Out(bn13_Data_Out),
		.Valid_Out(bn13_Valid_Out)
	);
	Relu_Core rl_kernel13(
		.Data_In(bn13_Data_Out),
		.Valid_In(bn13_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(rl13_Valid_Out)
	);
//////////KERNEL14//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111110110000001110010110000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111110100101001101110010000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110011110010000100111000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111100111011001001100101011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111110110011110001101000100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110110110111100000101001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111111000000100100011111110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111111000100011111011001101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110110110100001100100110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111111000000011100111011001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111111000101100001001101100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111011101100000111101000110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111110100000110101001100010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111110111011111111000011000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110101100101101100100111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111101101000110001001001111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111111010011001110111111100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111101101001101011100010000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111101001111000000100011100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111011110111000100000111111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110001001100011101011101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111110111101111110000111100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111101110110100111110001100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111101111100101110110110001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111101101000001010110110001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110100101100001000010111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111110111110011000111011100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110100011010111000101010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111111000000100101011111110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110000001110010110100111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111110111101010010010010000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111010000100110110010101010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b00111110000111111000010000101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b00111110100101011110111110110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111110001011111110110111000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b10111111001000010101001100111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111110010011100000011100000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111111001111010001101100101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b00111111011111111000110100111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b00111101100111110011101111100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111110100110101010111101011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b10111110010100110111001110000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111110100101011001111101011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111110110111001110110011101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b00111110101001010010111100011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b10111101011000100010100110110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b10111110000111011111010101010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b00111111000010011101101000011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111101100101010001001011101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111111000110110001001100110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111110010110000100010110010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b10111101101101100001011101011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111100111010011010101010010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b00111111010001011110001011001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111101101000110101100110000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b00111110101111010010000000110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111110001011111011111001010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b10111110001111110000000100111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b10111110110111110011110101011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111110110111011110010101011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b10111111000111000101011101111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b10111110010001101001101000101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111110010100110110111110001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b10111101101100110001000001111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel14_Valid_Out)
	);
	Adder_64input add_k14(
		.Data1(Data_Out_Kernel14[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel14[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel14[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel14[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel14[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel14[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel14[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel14[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel14[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel14[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel14[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel14[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel14[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel14[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel14[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel14[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel14[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel14[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel14[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel14[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel14[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel14[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel14[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel14[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel14[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel14[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel14[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel14[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel14[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel14[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel14[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel14[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel14[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel14[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel14[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel14[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel14[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel14[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel14[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel14[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel14[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel14[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel14[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel14[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel14[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel14[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel14[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel14[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel14[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel14[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel14[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel14[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel14[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel14[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel14[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel14[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel14[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel14[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel14[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel14[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel14[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel14[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel14[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel14[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel14),
		.Data_Out(add_k14_Data_Out),
		.Valid_Out(add_kernel14_Valid_Out)
	);
	Batch_Norm bn_kernel14(
		.Data_A(32'b00111111000000011010101011000111),
		.Data_B(32'b00111110001000101011100100111011),
		.Data_In(add_k14_Data_Out),
		.Valid_In(add_kernel14_Valid_Out),
		.Data_Out(bn14_Data_Out),
		.Valid_Out(bn14_Valid_Out)
	);
	Relu_Core rl_kernel14(
		.Data_In(bn14_Data_Out),
		.Valid_In(bn14_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(rl14_Valid_Out)
	);
//////////KERNEL15//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111110010101110011010010010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110101110010101101100001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111100011101101011000101001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110110000110110001000100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111110100110000110100011110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110001010111000010000001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111110001111010100000000010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111110011100001001000101011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111110111100100110100010011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111101000100000011001010101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111101100010001001110011100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111101001011000011100000110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111101110000101101000000001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111101101010111100110100111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110110101101100000001110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111101010101010111011100000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111111010110111010101010100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111101110101110111010001011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111110110000111011011001111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110000001100001000001011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111111001111001010110101000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111110001111001000000000010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111110011010001000100010010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111110100011100110110001101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111101101011011001001011001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111110000011101100001101001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111111000101101000011010010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111110000111000000010011101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111110110000110011101110001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110111000111100100110010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111110001100100111001101101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111101001101111101011101011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b00111101110111110011110011110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b00111101111110000010001111000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111111000001000101010110010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111101111101011110100101110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111101010101001001010101011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b00111110110110111100000000110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111111010110000011001001000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111101011101101011011110101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111101000111111001101111010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111111010100111010101010110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b00111110101111101001110001000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b00111110011111100001000001111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b00111110100000011100011101101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111101000101101011101111001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b10111111011011001110100100010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111110101010101100010001110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111110111101110101000010011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b00111110001110110101001010001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b10111101010000001011000010011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111110101010001010100110010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b00111111011111100010111111100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111110010111100111100001111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111101101000101110100110011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111110000100110010110101001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111110101110011000001000101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b10111110001101111000101111000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111101110101001111010011110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b00111111001010010111011110111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b10111110110101000010000001111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111110001011001001000101101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111110100101111001011010010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111101111111010011100111111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel15_Valid_Out)
	);
	Adder_64input add_k15(
		.Data1(Data_Out_Kernel15[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel15[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel15[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel15[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel15[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel15[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel15[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel15[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel15[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel15[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel15[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel15[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel15[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel15[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel15[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel15[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel15[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel15[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel15[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel15[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel15[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel15[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel15[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel15[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel15[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel15[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel15[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel15[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel15[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel15[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel15[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel15[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel15[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel15[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel15[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel15[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel15[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel15[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel15[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel15[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel15[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel15[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel15[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel15[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel15[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel15[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel15[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel15[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel15[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel15[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel15[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel15[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel15[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel15[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel15[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel15[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel15[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel15[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel15[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel15[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel15[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel15[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel15[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel15[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel15),
		.Data_Out(add_k15_Data_Out),
		.Valid_Out(add_kernel15_Valid_Out)
	);
	Batch_Norm bn_kernel15(
		.Data_A(32'b00111110110101000010011011111011),
		.Data_B(32'b00111101100000010001100100011100),
		.Data_In(add_k15_Data_Out),
		.Valid_In(add_kernel15_Valid_Out),
		.Data_Out(bn15_Data_Out),
		.Valid_Out(bn15_Valid_Out)
	);
	Relu_Core rl_kernel15(
		.Data_In(bn15_Data_Out),
		.Valid_In(bn15_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(rl15_Valid_Out)
	);
//////////KERNEL16//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111110001010000101110000000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111110111100111000111100101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111101010111100100000100001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110001001100100101100000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111110011011101011000110010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111101110011010001011101111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111110011100110011001000110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111111000101111000010000000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111110101000111100101001001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111111000101100001111000111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111110101110100110111111010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111101001100010011000101001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111111011001001000001010111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111111000000011001101001110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110101000011101010001111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111110100101100110001000111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111101011011010010001111010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111110000000111110010011100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111111000100011111011000010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110001110001101100000111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111111000110100010010101010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111110101111111001000101010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111110101010100100001110000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111110100110110100000001001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111110000001010011100000010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111101101110011111000011000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111111001001111011110000011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111111001000111110101001010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111101001011001001010010010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111110111110000110011000101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111110100010000001111110100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110110110101111111000011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b00111111001101000001100010111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111100111100101101011101110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111110111010100100101100000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111110000011000110111101000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111101100001011101000001000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111110110111010011010110000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b00111100111111001010100100011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111111001101011110001010101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111100101001010011011101001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111110111010011000100101010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111100001101000011011101110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b00111110010001100001101110000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b00111110010010001011001100000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b10111101110001010101011011001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b10111110110001010000000100011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b00111110110001110111100110111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111110010010011001011111111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111110001001101100001010111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111111000011010001001110010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111101100100001100010011010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111110011101001101001000100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111110011011110111010010000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111110010001100110000111100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b00111110010011100110101011101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111110100100010001101010110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111110100111001101111010010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111110111100000110010011000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b00111110101011110001110001011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111101111001010001001011100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111110011110000011001111101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b10111110000101100000110110110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b10111110110110111010111100000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel16_Valid_Out)
	);
	Adder_64input add_k16(
		.Data1(Data_Out_Kernel16[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel16[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel16[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel16[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel16[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel16[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel16[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel16[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel16[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel16[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel16[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel16[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel16[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel16[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel16[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel16[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel16[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel16[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel16[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel16[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel16[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel16[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel16[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel16[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel16[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel16[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel16[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel16[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel16[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel16[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel16[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel16[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel16[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel16[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel16[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel16[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel16[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel16[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel16[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel16[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel16[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel16[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel16[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel16[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel16[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel16[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel16[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel16[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel16[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel16[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel16[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel16[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel16[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel16[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel16[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel16[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel16[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel16[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel16[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel16[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel16[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel16[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel16[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel16[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel16),
		.Data_Out(add_k16_Data_Out),
		.Valid_Out(add_kernel16_Valid_Out)
	);
	Batch_Norm bn_kernel16(
		.Data_A(32'b00111110111000110110111011010110),
		.Data_B(32'b00111101110111110010001100101100),
		.Data_In(add_k16_Data_Out),
		.Valid_In(add_kernel16_Valid_Out),
		.Data_Out(bn16_Data_Out),
		.Valid_Out(bn16_Valid_Out)
	);
	Relu_Core rl_kernel16(
		.Data_In(bn16_Data_Out),
		.Valid_In(bn16_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(rl16_Valid_Out)
	);
//////////KERNEL17//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111110110101010111000110110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110110001011000110100100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111100110100000000111000101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111101000111110100100011010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111111000011110000000101011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111111001010010101100100101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111110011001110000001100010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111110111101100000011101010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111101100100000010011100111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111110001101110001010101010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110011110101101000101110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110000000001101010010111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111110010001000110011000101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111110100001011010100111000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110101010101000011111010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111110111000001000000010110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110011101101001100000111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110101100011010010110001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111110100000111011011100111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110000000001010101011100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110010101111101101111011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111110100011001110111110011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111100000100011011000110011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111110000011000111010100001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111101110101001000100001101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111101100001001110011011111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111111000110010010101111110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110101111011100111100010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111110101000001011110000110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110011111010110000110011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111110110110100110000000000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111111010001110000011101100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b00111110101100001100010011101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b00111110001110111000110000110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111110100001110010011100110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111111000101111011011011010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b10111111000111011100111011110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111110011111110111011111010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111110000110000010111101111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111111001001010000111111101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b10111110011110011110000010101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b10111101001110010101110110011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b00111110101000011010011000000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111111010111001101100001011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111111100000101001100110010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111110100101110101001100111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b10111101110001010101101101111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111110010011001011011111111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111011111111000101101110010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b00111110010111100011011101101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b10111110111000100100111101100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b10111101101010000010001001111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b00111110001010100000111001110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b00111101100101111100111000101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111110100010110001011110101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b00111110011000101111010001110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b10111111001110001111100011110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111110100101011101011011100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b10111110001111101111000101111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b00111110110010110111010111111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111100110010011000100001111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b10111101010101111000111011111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111110110010101101010110000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b10111110011101110101111001011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel17_Valid_Out)
	);
	Adder_64input add_k17(
		.Data1(Data_Out_Kernel17[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel17[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel17[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel17[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel17[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel17[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel17[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel17[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel17[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel17[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel17[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel17[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel17[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel17[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel17[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel17[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel17[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel17[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel17[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel17[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel17[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel17[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel17[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel17[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel17[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel17[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel17[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel17[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel17[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel17[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel17[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel17[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel17[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel17[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel17[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel17[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel17[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel17[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel17[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel17[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel17[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel17[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel17[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel17[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel17[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel17[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel17[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel17[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel17[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel17[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel17[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel17[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel17[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel17[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel17[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel17[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel17[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel17[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel17[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel17[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel17[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel17[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel17[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel17[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel17),
		.Data_Out(add_k17_Data_Out),
		.Valid_Out(add_kernel17_Valid_Out)
	);
	Batch_Norm bn_kernel17(
		.Data_A(32'b00111110111100110000010100101001),
		.Data_B(32'b00111111001100000010110111101100),
		.Data_In(add_k17_Data_Out),
		.Valid_In(add_kernel17_Valid_Out),
		.Data_Out(bn17_Data_Out),
		.Valid_Out(bn17_Valid_Out)
	);
	Relu_Core rl_kernel17(
		.Data_In(bn17_Data_Out),
		.Valid_In(bn17_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(rl17_Valid_Out)
	);
//////////KERNEL18//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111101100001010011101111111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111101110110100010110011000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111100110100011011010110110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111100110110000010010110011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111110101011111011110011101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111110011001010011101010100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111110000010110100111101011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111101100010011000100111001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110111010100011111001110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111111011001110000011100100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111111000010111100100110110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111111001001001111010111100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111110000001001010101001001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111110100110100010010100110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111101111111010010001100111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111110111000111011011100011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111110100001101111001011100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111010110010011001000011111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110101010001001100111110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111110100000011111001000010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111101000111000011000010010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111100011111111010011101111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111111001001010011100011000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111101100000101110011110100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111110101001000001101011111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110000101010001110111011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110100110110001010111011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111101110000100011000001100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111110001011101010100111100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110111011100101110100111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111110110011111100110001100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111111000000001001101101111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111110000101110010011011110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111100101010011111011100000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111111000110101011110000000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111110110000111001100110111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111111100110001100010101001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111110101111001111110101000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111101110100011011011000100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b00111111000000011000011100111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111101110001111100010110010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b10111101100110001101111101001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111110101100110011000111101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b00111110111101010001101011110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111110101100010100110111101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111110011010011110010000011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b10111110101001010000100100100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111110100001101101010100101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b00111110000001100000000110101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111110101111110100010010010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b10111101110000011011110101001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111110001001111001001111100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b00111101101011101000101001010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111110100111110110111011011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111110100001000001100000111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111110011010101111110011100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111110101000001001001101101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111111011111110010111010011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111110011000100001011111101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111110000101010101001000101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b10111011011011110100001010011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111110111110100010101100101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b10111110100000000001000000000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111110011101000011111100011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel18_Valid_Out)
	);
	Adder_64input add_k18(
		.Data1(Data_Out_Kernel18[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel18[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel18[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel18[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel18[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel18[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel18[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel18[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel18[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel18[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel18[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel18[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel18[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel18[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel18[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel18[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel18[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel18[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel18[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel18[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel18[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel18[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel18[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel18[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel18[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel18[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel18[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel18[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel18[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel18[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel18[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel18[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel18[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel18[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel18[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel18[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel18[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel18[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel18[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel18[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel18[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel18[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel18[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel18[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel18[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel18[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel18[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel18[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel18[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel18[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel18[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel18[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel18[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel18[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel18[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel18[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel18[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel18[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel18[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel18[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel18[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel18[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel18[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel18[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel18),
		.Data_Out(add_k18_Data_Out),
		.Valid_Out(add_kernel18_Valid_Out)
	);
	Batch_Norm bn_kernel18(
		.Data_A(32'b00111110110101000000111111100011),
		.Data_B(32'b00111111100001011110000100010010),
		.Data_In(add_k18_Data_Out),
		.Valid_In(add_kernel18_Valid_Out),
		.Data_Out(bn18_Data_Out),
		.Valid_Out(bn18_Valid_Out)
	);
	Relu_Core rl_kernel18(
		.Data_In(bn18_Data_Out),
		.Valid_In(bn18_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(rl18_Valid_Out)
	);
//////////KERNEL19//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110001010101011101010000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110010100100011010110100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110111011011111001011000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111111000000001100110110110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111110110001010011111000011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110110010111010110101001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111111000001000001000101000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111110000001111111001101000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110101101011111110100101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111110100101101101110100000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110100011001010101100110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111101100001110010100011001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111101111001110011011111011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111110000110111000101011110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110100110000100110000100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111011101010011000001011010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111101101110101010111001010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110101111000101000101000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110001001101111001011100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110110001101000010000101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110011101110101011101010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111101101110110110101110101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111110101011000110001111011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111101101011101000010110010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111101110010010100111000110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111101101110010101001010110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111101011011111100110011111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111101101110010010001110100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111111000011001101100101100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110001000001110011010001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111101111111111010110010010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110010010011000101010100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b00111111100100110010011001000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111110110100010000010101111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111110101001111111110111011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111111001110011101110011001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111110110001010000110001011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111110111011111000011110110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b00111101111000011010100001000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b00111111000110010100011011111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111111000011001101110000100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b10111110101011100011011000101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111110111110000000001001111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b00111101111010111011011011111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111110100000110101011111000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b10111110101100111111000011101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111110000101010100000110010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b00111110101001100011011001010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111110111110100000000101100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b00111101101101011111110010111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b10111110111001001001001001100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b10111111000111000111111010000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b00111100101110001010011011000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b00111111001011111010110011100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111110111110001110000100110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b00111110000110100000101001010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b10111110011010111001011010100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111111000001101111010001100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b10111101011111110111111011100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111101010110011100011110110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111110101110011111110110111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111110010000101010000110010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b10111101010000111110100000010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b10111111000011011011001010000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel19_Valid_Out)
	);
	Adder_64input add_k19(
		.Data1(Data_Out_Kernel19[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel19[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel19[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel19[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel19[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel19[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel19[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel19[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel19[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel19[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel19[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel19[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel19[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel19[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel19[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel19[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel19[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel19[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel19[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel19[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel19[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel19[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel19[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel19[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel19[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel19[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel19[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel19[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel19[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel19[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel19[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel19[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel19[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel19[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel19[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel19[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel19[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel19[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel19[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel19[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel19[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel19[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel19[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel19[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel19[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel19[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel19[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel19[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel19[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel19[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel19[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel19[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel19[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel19[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel19[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel19[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel19[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel19[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel19[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel19[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel19[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel19[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel19[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel19[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel19),
		.Data_Out(add_k19_Data_Out),
		.Valid_Out(add_kernel19_Valid_Out)
	);
	Batch_Norm bn_kernel19(
		.Data_A(32'b00111110111100000011000011110000),
		.Data_B(32'b00111111001001101100011110111101),
		.Data_In(add_k19_Data_Out),
		.Valid_In(add_kernel19_Valid_Out),
		.Data_Out(bn19_Data_Out),
		.Valid_Out(bn19_Valid_Out)
	);
	Relu_Core rl_kernel19(
		.Data_In(bn19_Data_Out),
		.Valid_In(bn19_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(rl19_Valid_Out)
	);
//////////KERNEL20//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110101001110000000010111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111111000101011010000100111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110100000000010111010000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111111000111001011100101101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111110010110100000001010001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111100110110011011000100010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111101111100010110110011100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111110100101011010100010101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110101010010100000111010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111101100101000111000101001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111111010011101000100101101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111101110101111101100001111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110000010100000110111000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111111001000000010100010101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111111000010001101010100000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111110011010010101110011010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110000010110011001111111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111111000001011001110100010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111100010100101000101000110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110111011110001101101010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110100110111010110000000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111110100110100111001010111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111111001010010101001001001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111110101000110011110100101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111101111011111000011001110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110111101001110110100010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111101101101101111100101100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111111001110011010000010110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111100101010110110110010101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111110011011001100111111111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111110001110001000000010000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111101011000001001010100010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b00111101111100011101001000000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b00111110110110001101111010000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111101100101010100000001100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b10111110100101001111011011101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b10111110110010010101111111101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b00111110100010110101101111010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b00111110101101010110110100100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111101101011000100110000100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111110011110010010101101111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111110101101111100011101110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111110000001001110001100101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b00111111000111111010011010101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111110100110011111001001110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b10111110110111111110000010010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111110110101000010000111010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111111000010101011101111011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b00111110110110101111111010001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111111100011011010011010010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111110001011110011001100100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b10111101111011001010100011010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111101011010001001101010110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111111010100100101110001010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b10111011110001101110010100000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b00111110011001000100100000100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b10111101011111100010000100010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b10111101101011110100101101101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111100101101011010101010101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111111001000111100111000100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b10111110111011101000000111001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b10111110110110011010001111001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111110010011110101111010010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b10111110001111011000001110001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel20_Valid_Out)
	);
	Adder_64input add_k20(
		.Data1(Data_Out_Kernel20[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel20[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel20[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel20[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel20[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel20[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel20[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel20[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel20[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel20[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel20[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel20[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel20[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel20[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel20[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel20[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel20[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel20[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel20[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel20[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel20[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel20[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel20[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel20[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel20[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel20[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel20[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel20[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel20[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel20[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel20[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel20[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel20[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel20[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel20[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel20[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel20[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel20[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel20[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel20[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel20[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel20[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel20[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel20[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel20[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel20[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel20[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel20[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel20[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel20[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel20[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel20[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel20[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel20[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel20[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel20[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel20[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel20[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel20[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel20[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel20[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel20[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel20[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel20[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel20),
		.Data_Out(add_k20_Data_Out),
		.Valid_Out(add_kernel20_Valid_Out)
	);
	Batch_Norm bn_kernel20(
		.Data_A(32'b00111110110100011101010011111000),
		.Data_B(32'b00111111011010000001011011101011),
		.Data_In(add_k20_Data_Out),
		.Valid_In(add_kernel20_Valid_Out),
		.Data_Out(bn20_Data_Out),
		.Valid_Out(bn20_Valid_Out)
	);
	Relu_Core rl_kernel20(
		.Data_In(bn20_Data_Out),
		.Valid_In(bn20_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(rl20_Valid_Out)
	);
//////////KERNEL21//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110111111010000110101011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111101000110011110010000100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111100111010010100100100010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111111000000001110111110001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111111010010010011111010101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111111011110101110000101001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111100101010001110100111000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111111000000010010111100100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111111010000110010001011110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111110001001010011011000000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111110100011010101010101110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111110011110110101000101100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111110010000111111101111011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111100101110011001110111101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111101101000011111100011100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111101011000000011100001001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110110100100000000111101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110100001111011010011100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111100100101010010010100100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110110001110100110010110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111101110001110010110011101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111110001000010000111010010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111101110100011101101001011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111101110110100100110110000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111110110001100011100101111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110100111111011001101111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111100110010001010100101010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110010011101011111011110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111101111000010001110000100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111110101010101010000101100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111110111000110110110110100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111011011101011011100001111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b00111110100110011001101001010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111111000010000001010001100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111110001011010010100001001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111111010110100011001110111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111111000001010110000011000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b00111110110001000111011100010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111110101111001010011001010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111111000110011001110111011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b10111110100001101000100001111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111101111000011101110100111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111110100000011011100010011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b00111101010101110101111111010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b00111100101101011001101100001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111101000011001101010001110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b10111111000100000011010001001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111101000011100001100010011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111110111011001010110011010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b00111101010001001110000111110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111110001110001000010000000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111111001011000000110101110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b00111110100100101111011011101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b00111110011001001000100110010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111101011011100001011000011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111110010110000000101110011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111101100101000100011110000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111100001001010000100010101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b10111111011011000110100110001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111101001011101100011101010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111101111001111000111111110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111101010111101100001011101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b10111101011110101011111101111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b10111110011010001101011010101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel21_Valid_Out)
	);
	Adder_64input add_k21(
		.Data1(Data_Out_Kernel21[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel21[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel21[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel21[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel21[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel21[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel21[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel21[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel21[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel21[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel21[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel21[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel21[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel21[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel21[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel21[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel21[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel21[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel21[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel21[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel21[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel21[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel21[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel21[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel21[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel21[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel21[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel21[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel21[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel21[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel21[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel21[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel21[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel21[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel21[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel21[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel21[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel21[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel21[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel21[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel21[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel21[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel21[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel21[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel21[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel21[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel21[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel21[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel21[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel21[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel21[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel21[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel21[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel21[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel21[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel21[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel21[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel21[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel21[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel21[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel21[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel21[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel21[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel21[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel21),
		.Data_Out(add_k21_Data_Out),
		.Valid_Out(add_kernel21_Valid_Out)
	);
	Batch_Norm bn_kernel21(
		.Data_A(32'b00111110111000000000110000001001),
		.Data_B(32'b00111110111110011110111111001010),
		.Data_In(add_k21_Data_Out),
		.Valid_In(add_kernel21_Valid_Out),
		.Data_Out(bn21_Data_Out),
		.Valid_Out(bn21_Valid_Out)
	);
	Relu_Core rl_kernel21(
		.Data_In(bn21_Data_Out),
		.Valid_In(bn21_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(rl21_Valid_Out)
	);
//////////KERNEL22//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110100010011000111110011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110001001110000000111101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110110110011111010001011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110010100011001000111101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111110101011001010111111101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111110000101010111110100100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111101110110010100110000000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111110111000101110110111001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110111001111100011111011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110010110100111110110011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111110000100101111110010101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111111001010100001100011000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111010110110111010110011100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111110000010111100100100101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110100000001010101100001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111110110000010111111110110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111111000101000110000101110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111110100100001001000010010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110010101000101110101110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111111010011000010001100011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110101010111010100011101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111111001010010000111000101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111110100010001000000000001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111111010000100000111111011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111100110111010100100111000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111011110010011110110100000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111101111100100100101111011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111111000011011110011101100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111110111100111100001101110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110110000101100001100101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111110001110000000010000100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111101111011110110100110100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b00111110110110101111111001101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111110000001011010111101100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111110010110000000110000010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b10111110001110100001101011100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111110010001100100001100010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111110001110010100010111001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111101101100101110111100101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111101101110101101011110000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111111010011100110111111001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b10111111011001001100111011011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b00111101111101101101010011010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b00111101101110010100100111101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111110001001100100110110010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111101100110101010111010100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111110111000101001101000100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b00111110011101011001010010100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111100110101010101110101010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111110100110001001100100010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b10111110001110000011110010101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111110111001001111001000111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b00111111001111011001101011110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111110101010110000001001001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111110101100000110010000100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b00111110111110111101010000001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111110111010110001001101101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111101101100000110010011010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b10111110100011000000011001101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b00111110111011000100011111111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111110001001010110000111100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111110010111101101101100000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111110100100101011001110001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b10111111000010000101001001001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel22_Valid_Out)
	);
	Adder_64input add_k22(
		.Data1(Data_Out_Kernel22[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel22[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel22[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel22[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel22[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel22[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel22[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel22[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel22[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel22[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel22[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel22[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel22[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel22[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel22[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel22[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel22[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel22[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel22[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel22[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel22[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel22[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel22[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel22[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel22[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel22[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel22[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel22[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel22[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel22[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel22[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel22[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel22[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel22[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel22[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel22[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel22[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel22[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel22[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel22[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel22[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel22[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel22[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel22[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel22[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel22[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel22[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel22[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel22[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel22[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel22[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel22[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel22[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel22[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel22[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel22[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel22[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel22[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel22[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel22[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel22[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel22[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel22[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel22[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel22),
		.Data_Out(add_k22_Data_Out),
		.Valid_Out(add_kernel22_Valid_Out)
	);
	Batch_Norm bn_kernel22(
		.Data_A(32'b00111110110010011111010010010100),
		.Data_B(32'b00111111010010101010011110111011),
		.Data_In(add_k22_Data_Out),
		.Valid_In(add_kernel22_Valid_Out),
		.Data_Out(bn22_Data_Out),
		.Valid_Out(bn22_Valid_Out)
	);
	Relu_Core rl_kernel22(
		.Data_In(bn22_Data_Out),
		.Valid_In(bn22_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(rl22_Valid_Out)
	);
//////////KERNEL23//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111101110110001000101111010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110011011000000011000110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111111010110100111100110110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110101000000000010000100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111110000000110011000011111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111110111011101010110101010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111111000001101000000011100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111101000100011101100001011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111110010100111011001110111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111110010100110110101000111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111110100001010101111101001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110001111110100000010110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110001011111001101011110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111110000101101100010100011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110000110011001111011111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111110010110101110101111111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110011000001000110101010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111101110100010010001100110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111111000000111111010011010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111100101111100001110011100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111101101011001011001001100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111110110101111011011011010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111101110111100100111010010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111110011101101110000000011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111110000010111111110111111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110101000110010010000001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111110100101110110100110101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111110010110110111000000100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111110100101110111001011011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111110101010111011000001011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111111000000010000001110110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111111010001111010101011110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b00111100101111101110111000011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b00111110110011100110111001101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111111001111101000001101110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111110101011100110010011001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b10111110101101110100000010011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b00111110100011111100011100001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b00111110101101100010010110110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111110001101011101101011101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b10111110000011000000110100011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111101011100110111001000011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b00111111000001110001001010100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111110100101110100010001011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111111001110000010110100011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b10111110100100101111101000100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b10111101010011110111011100100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111110111111011000000101011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b00111101011011000000001001011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111101100001101010001100101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b10111110110100110100011100010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111101101100001001100011101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b00111110111110000111000110100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111110110110000010101101010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111101111111101001010111110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111110101100011110010000011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b10111111010001101000010101110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111110100101010000110111111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b10111110111111000100011000101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b00111110001011100010001111000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b10111101110010111110011000101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b10111111000101110110000000001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b10111101010000110011101110110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111111000001100101011101001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel23_Valid_Out)
	);
	Adder_64input add_k23(
		.Data1(Data_Out_Kernel23[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel23[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel23[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel23[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel23[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel23[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel23[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel23[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel23[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel23[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel23[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel23[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel23[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel23[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel23[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel23[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel23[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel23[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel23[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel23[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel23[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel23[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel23[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel23[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel23[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel23[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel23[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel23[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel23[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel23[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel23[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel23[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel23[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel23[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel23[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel23[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel23[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel23[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel23[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel23[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel23[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel23[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel23[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel23[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel23[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel23[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel23[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel23[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel23[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel23[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel23[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel23[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel23[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel23[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel23[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel23[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel23[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel23[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel23[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel23[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel23[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel23[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel23[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel23[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel23),
		.Data_Out(add_k23_Data_Out),
		.Valid_Out(add_kernel23_Valid_Out)
	);
	Batch_Norm bn_kernel23(
		.Data_A(32'b00111111000000100011010111100001),
		.Data_B(32'b00111111001000000001000101100111),
		.Data_In(add_k23_Data_Out),
		.Valid_In(add_kernel23_Valid_Out),
		.Data_Out(bn23_Data_Out),
		.Valid_Out(bn23_Valid_Out)
	);
	Relu_Core rl_kernel23(
		.Data_In(bn23_Data_Out),
		.Valid_In(bn23_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(rl23_Valid_Out)
	);
//////////KERNEL24//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110000000101001101101100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111110110110010101010101111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110100110000101100111110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110011011100101100000000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111110100001011001011111101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111110010111001010110110000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111110011111001010010010100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111110100110111100110011000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111111010011100101001011000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110111110010000011101101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111110001010100110110110100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110011100000110101000010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111110100010111010001001101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111100111011001110010101110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111101110111111110100000101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111100101000111101101110101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111110111111000101001110010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111111000110011011010001110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110100101101111010011001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111110010110011110110110000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110001110100111011000111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111110110110101111011011011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111110101001100101111101000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111110001101000010110100000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111110000010100110100001011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110111101101100110001101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110001001101000100010000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111101111011010010010110111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111111001110110110100000101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111101101001101101010010011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111110001101001000100100010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111110001010100100111011111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b00111110000111100000001111110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b00111111000110111100100000000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111110000111010000111110101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b10111110101000101110101100100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b10111110011100000101100111100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111110010000100101110111000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b00111111000001001101010110010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b00111110111100010111100011011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b10111111000101011110000010011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b10111110101011111010100100101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b00111111010100001001110001011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b00111110111010011001001101100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b00111100100011001010010001110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b10111101101000010100110101101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111110101111111100111101010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b00111011111100000001101001110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b00111101111001100100100101110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111101101111100011001000010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b10111110101001100001011000100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b10111110111010001001010010101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b00111101011010110010100110000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111110101111011101010101011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111110000110101011000011010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111111001110101001001000110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111101010010111010110101011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111101010110000111110010111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b10111110000110000001010010101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111111000100100001001100000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111110110111010000100100111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111110111011001001101001101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b10111111001111110110001001110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b10111101001000111100010110011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel24_Valid_Out)
	);
	Adder_64input add_k24(
		.Data1(Data_Out_Kernel24[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel24[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel24[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel24[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel24[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel24[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel24[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel24[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel24[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel24[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel24[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel24[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel24[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel24[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel24[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel24[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel24[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel24[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel24[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel24[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel24[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel24[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel24[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel24[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel24[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel24[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel24[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel24[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel24[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel24[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel24[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel24[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel24[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel24[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel24[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel24[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel24[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel24[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel24[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel24[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel24[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel24[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel24[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel24[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel24[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel24[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel24[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel24[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel24[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel24[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel24[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel24[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel24[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel24[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel24[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel24[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel24[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel24[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel24[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel24[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel24[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel24[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel24[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel24[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel24),
		.Data_Out(add_k24_Data_Out),
		.Valid_Out(add_kernel24_Valid_Out)
	);
	Batch_Norm bn_kernel24(
		.Data_A(32'b00111110111000110100101110100001),
		.Data_B(32'b00111101001011011001110101110101),
		.Data_In(add_k24_Data_Out),
		.Valid_In(add_kernel24_Valid_Out),
		.Data_Out(bn24_Data_Out),
		.Valid_Out(bn24_Valid_Out)
	);
	Relu_Core rl_kernel24(
		.Data_In(bn24_Data_Out),
		.Valid_In(bn24_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(rl24_Valid_Out)
	);
//////////KERNEL25//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110010001011110011101010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111110001111100011001001101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110110000000011110000101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110101001001010101010110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111110010000100110010000011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110011101111111010001000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111111000000101110001010111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111101100010110100010010111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111110110000010111001011011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110101011001110010101001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111110101101010010010000111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111110110000010001101001111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111110010101111100000101001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111110011000011011001111010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110101101000101100101010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111101110010110110000010011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110101111001011010100110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111111001011010011100001101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111101111100000000001111011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111111010100011110001110001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111101010100011000100000101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111110000010001111001001100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111101000110010011001000011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111101001101110001110110111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111101101010101110001011000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110000100111110110011010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111111000011111001001110111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110111101101000110000110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111101011010011011010011111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111110101000110111011111100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111110000000001000110110010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110111010000000110000000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111110110001111101011100010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111110100011000011001001011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111111000010100100100111100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111101110110110011101110011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b10111100101111001101110110000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111110101010011101110000010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b00111110100000001000011111001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b00111110101000010101111110011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111011111000110111001011101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b10111101110010110100000000101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111110101101010100001111011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b00111111000011111011011010100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b00111110000010101000100001000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111100101000011010100011100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111110010011011011101000000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b00111110000000100100010111011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b00111101000111101011011011101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b00111101011000001011111001110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b10111110101011010110111100000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111111001011001100001011111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111111000110100010001011011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b00111110100010001101001010110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111111001011001010010011010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b00111110110111010101001101101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111111001001011100001111111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b10111100010111111011100110110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b10111110011101111101101110100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111110110111011001010011011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b10111111000000101011001101100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111110111011110111100110010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111111000000101000110101100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111101111110100000000100101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel25_Valid_Out)
	);
	Adder_64input add_k25(
		.Data1(Data_Out_Kernel25[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel25[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel25[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel25[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel25[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel25[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel25[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel25[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel25[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel25[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel25[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel25[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel25[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel25[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel25[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel25[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel25[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel25[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel25[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel25[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel25[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel25[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel25[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel25[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel25[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel25[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel25[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel25[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel25[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel25[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel25[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel25[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel25[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel25[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel25[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel25[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel25[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel25[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel25[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel25[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel25[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel25[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel25[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel25[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel25[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel25[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel25[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel25[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel25[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel25[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel25[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel25[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel25[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel25[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel25[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel25[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel25[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel25[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel25[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel25[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel25[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel25[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel25[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel25[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel25),
		.Data_Out(add_k25_Data_Out),
		.Valid_Out(add_kernel25_Valid_Out)
	);
	Batch_Norm bn_kernel25(
		.Data_A(32'b00111111000001000110000010101000),
		.Data_B(32'b00111110101110000111001011100100),
		.Data_In(add_k25_Data_Out),
		.Valid_In(add_kernel25_Valid_Out),
		.Data_Out(bn25_Data_Out),
		.Valid_Out(bn25_Valid_Out)
	);
	Relu_Core rl_kernel25(
		.Data_In(bn25_Data_Out),
		.Valid_In(bn25_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(rl25_Valid_Out)
	);
//////////KERNEL26//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111110111011000001000111101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111101000111001000010101110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110011111001001011111101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110100111111000011101101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111100100100011011101011110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111110110010000011100011011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111110111001101101000110111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111110010011010111110001011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111110100000010101010100000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110011100011000100000011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110100111011110100000010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111111000011110010110111100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110100101100101111101000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111110111101100000110000101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111101100101001011011011011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111101001010001000110010101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111110101100101001000010110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111110100101100000101011001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111101100110010110011001111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110101110011000100101010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110011010110101010001010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111110100111000111111111010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111101100100001101010100011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111110001111011000101101001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111110101011010100001010010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111111010110111101101000100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111110110000100011011010100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110101011100111001000110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111110110111010011010100101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110001101110101101101101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111101101011100110100101000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111110100110110011000001100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b00111110100010111001111110110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b00111101111111111111101110111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111110100011110101111011010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b10111100100011000001001110110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111110110001110110100110010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b00111111000010111001011010011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111110001010010100010110000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b00111101101111100011110010100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b10111110010110010100110011101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111111001011100110010000100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111110001110010001101100011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b00111101000100111100001110000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111110000010010011001011100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111110111011110001111111110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b10111101111001110101010000010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b00111110100100000010011001100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111101110001000101001000101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111110100010000000010001111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111101000101011000000000101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b10111111000010001010100010000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111101110100001110100001001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111101101000111100101111101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b10111111000110000111001101010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b00111110000111001111111000101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111111000001101010110100010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111100111010011110001010111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b10111111000111101000000001010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b00111101000110100110100100011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111110110100110010111110011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111111000100111000101001010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b10111111011010010000011101000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111111000001100000100010110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel26_Valid_Out)
	);
	Adder_64input add_k26(
		.Data1(Data_Out_Kernel26[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel26[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel26[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel26[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel26[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel26[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel26[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel26[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel26[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel26[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel26[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel26[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel26[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel26[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel26[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel26[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel26[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel26[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel26[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel26[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel26[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel26[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel26[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel26[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel26[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel26[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel26[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel26[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel26[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel26[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel26[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel26[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel26[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel26[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel26[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel26[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel26[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel26[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel26[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel26[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel26[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel26[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel26[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel26[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel26[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel26[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel26[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel26[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel26[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel26[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel26[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel26[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel26[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel26[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel26[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel26[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel26[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel26[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel26[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel26[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel26[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel26[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel26[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel26[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel26),
		.Data_Out(add_k26_Data_Out),
		.Valid_Out(add_kernel26_Valid_Out)
	);
	Batch_Norm bn_kernel26(
		.Data_A(32'b00111110111100001010011100101010),
		.Data_B(32'b00111110100011101100110001011001),
		.Data_In(add_k26_Data_Out),
		.Valid_In(add_kernel26_Valid_Out),
		.Data_Out(bn26_Data_Out),
		.Valid_Out(bn26_Valid_Out)
	);
	Relu_Core rl_kernel26(
		.Data_In(bn26_Data_Out),
		.Valid_In(bn26_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(rl26_Valid_Out)
	);
//////////KERNEL27//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110000111110010101110101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111111000000111101111101001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110011011001010100001010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111101011100000011011011110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111110010111110010100111010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111110000011001011010010100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111111000111101110011110011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111110101010000111101111001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111101111101101111110011110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111111001010100101000100000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111111001001000000010110100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110110011001010111011001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110100011011011101101101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111110011010101101111000111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111100111000110100100010010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111110100010011011111101000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111111010000111011111000101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111111000101001110100111110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111101111010001010001001111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111101111001000111010000100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110111100111010010011000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111100101101110111111010000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110100001000001100110100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111101001001111111100001001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111101111101100100001111111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111111000010110001101000000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111110111101010110110010000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111101011001000111110110011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111011101110001010010000101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111110001000101110100100100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111111000011001110101111010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111101011111011010000100101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111110011011000001110100110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111111001000000011000101100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111101100001000011100101111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111110100110111111000010001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111100010100001000000011110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111110011111001100100000000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111101001110001011111111111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111110010010100111001011001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111110100011001111110011011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111110111101000110011100000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111110010000011100110101011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111111000000001000111000000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111111000011100110110001111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b10111100110001100100000000110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111111001110000001101011000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111110110111110001110010011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b00111110000101101100110011100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b00111110000110000101011101100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111011110110011001100000010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b10111110101110000000101111101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111111000011000111011001011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111110111101110110000111010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111111000101101100011100111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b00111110101011001100110100010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b10111011101101000000000011110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b10111101111110011010101110100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b10111111001001110000011101111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b00111110011110101101110110101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b10111110101101100101100011101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111110101000111100110001010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b10111111000011101011111110001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111110010111101010000011001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel27_Valid_Out)
	);
	Adder_64input add_k27(
		.Data1(Data_Out_Kernel27[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel27[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel27[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel27[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel27[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel27[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel27[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel27[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel27[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel27[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel27[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel27[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel27[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel27[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel27[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel27[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel27[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel27[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel27[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel27[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel27[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel27[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel27[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel27[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel27[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel27[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel27[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel27[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel27[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel27[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel27[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel27[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel27[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel27[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel27[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel27[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel27[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel27[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel27[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel27[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel27[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel27[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel27[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel27[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel27[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel27[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel27[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel27[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel27[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel27[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel27[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel27[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel27[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel27[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel27[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel27[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel27[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel27[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel27[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel27[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel27[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel27[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel27[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel27[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel27),
		.Data_Out(add_k27_Data_Out),
		.Valid_Out(add_kernel27_Valid_Out)
	);
	Batch_Norm bn_kernel27(
		.Data_A(32'b00111110110111100000001100101011),
		.Data_B(32'b00111111001100101010001001101100),
		.Data_In(add_k27_Data_Out),
		.Valid_In(add_kernel27_Valid_Out),
		.Data_Out(bn27_Data_Out),
		.Valid_Out(bn27_Valid_Out)
	);
	Relu_Core rl_kernel27(
		.Data_In(bn27_Data_Out),
		.Valid_In(bn27_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(rl27_Valid_Out)
	);
//////////KERNEL28//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111100101001011110010010101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110111110000001010101110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111111000100111111101101000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110011100111111110011010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111110110111110100010011110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110010101010001000111110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111110100100000010101000101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111101001111100010011000011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111101110000010101101100000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111110111100011010101101000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111110011000011100111011010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111101000001101011000001101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111110000100101011011111101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111110100100001110101110000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110101000100000000111000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111110101100000010011100100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111110110100100000111011011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111111000001001010010111001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111111000101100011100010001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111110100110101001011100110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110100101100011001110000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111101101010011001000000111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111111000110000000111011010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111101110010101011101101010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111110110110001101101000010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110100100100100100111001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110111011001010000011101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111111011011101100110001101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111110101111100010100000110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110101011110110110110100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111111001010111000110100011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111111010000101101001111100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b00111110111100001100000101000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b00111110001011100011010000011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111101100101111010100110101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111110101001100101011010100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b10111100111100010110111011110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111111001010000111010000000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111111000011100101100000111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b00111101100100011001100011100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b10111110001100011110001000110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b10111110001001110100001101101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111110101011110001010010101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b00111111000110011000001111010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b00111111010111111101100000000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b10111110010010100001001000001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111110110001111100111101100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b00111110110101110001001101010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b00111110011010001001110001000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b00111101000110010100111010000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b10111110000110110100011111110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b10111110000110101110000111110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b00111110011100101110000000011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b00111110101101100011111101111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111101011010100100110011010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111100101100000111010010000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b10111110101011100000101001001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b10111110101101100010001001001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b10111110111010010101110110010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b00111110010111101110000101001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b10111110101001000111111010100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111110110000011101111100101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111110010111000101010110100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111110100010010011001001010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel28_Valid_Out)
	);
	Adder_64input add_k28(
		.Data1(Data_Out_Kernel28[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel28[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel28[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel28[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel28[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel28[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel28[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel28[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel28[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel28[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel28[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel28[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel28[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel28[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel28[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel28[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel28[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel28[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel28[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel28[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel28[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel28[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel28[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel28[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel28[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel28[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel28[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel28[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel28[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel28[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel28[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel28[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel28[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel28[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel28[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel28[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel28[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel28[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel28[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel28[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel28[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel28[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel28[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel28[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel28[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel28[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel28[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel28[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel28[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel28[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel28[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel28[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel28[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel28[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel28[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel28[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel28[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel28[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel28[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel28[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel28[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel28[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel28[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel28[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel28),
		.Data_Out(add_k28_Data_Out),
		.Valid_Out(add_kernel28_Valid_Out)
	);
	Batch_Norm bn_kernel28(
		.Data_A(32'b00111110110010111100111011000000),
		.Data_B(32'b00111111001010110001110001011100),
		.Data_In(add_k28_Data_Out),
		.Valid_In(add_kernel28_Valid_Out),
		.Data_Out(bn28_Data_Out),
		.Valid_Out(bn28_Valid_Out)
	);
	Relu_Core rl_kernel28(
		.Data_In(bn28_Data_Out),
		.Valid_In(bn28_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(rl28_Valid_Out)
	);
//////////KERNEL29//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110101010110000010110101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111101100000011101101110110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111111011000101101110101010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110100011110001000101001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111100101001001100101001110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111101000111011001110001110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111111000011011110101100010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111110010000010001110110100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110010101011010010010011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110101011001101111110110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110101110011101111010101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111110010011101011100000010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110100011010011010110011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111110000011110001000101010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111111100001101110100101101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111101111100100100010001111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110000101001000011111010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111110000111010011011111001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111110100110111100111100011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111110010010100111011110001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110111101101100001110111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111110100110000000001001110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111111000101000011110001011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111101100000000101101101100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111110111100001000011001001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111101101000000011110010011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111111000101100011001011110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111111001110100000101000110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111110100100110000110001110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111110010111001001100011111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111110101010001111101011110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111110000111010100111111010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111110100111000000110000011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111111000110001101100100110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111110111101111001001000001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b10111110011101110000101100001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b10111101110101110101010011101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111110010010010011100000001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b00111110001110011100001010001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111111001010000100011000010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b10111101010111111111001101000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b10111110110010100000110101101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b00111111001110011100110101100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111110000111000100000101100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111110100001011011000001110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111110110001111100110110001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b10111101111110101000011010010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111110101001100000101011001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b00111111100001001111101001100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111100101001110010000011011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111110011011001001110110111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b10111110100110001011000101100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b00111110101010111000110100010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b00111101000100001011100000111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111110011001101110101001110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b00111100101101000110110010000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b10111111000111000011001001110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111110100101011101101111000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b10111111001001001010101111001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111110000111111010101000111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111110000010011110111100101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b10111110000100100001111010000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111101101111001110111100011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111110001110111010110110100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel29_Valid_Out)
	);
	Adder_64input add_k29(
		.Data1(Data_Out_Kernel29[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel29[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel29[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel29[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel29[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel29[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel29[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel29[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel29[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel29[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel29[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel29[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel29[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel29[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel29[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel29[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel29[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel29[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel29[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel29[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel29[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel29[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel29[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel29[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel29[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel29[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel29[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel29[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel29[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel29[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel29[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel29[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel29[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel29[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel29[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel29[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel29[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel29[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel29[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel29[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel29[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel29[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel29[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel29[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel29[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel29[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel29[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel29[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel29[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel29[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel29[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel29[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel29[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel29[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel29[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel29[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel29[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel29[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel29[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel29[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel29[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel29[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel29[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel29[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel29),
		.Data_Out(add_k29_Data_Out),
		.Valid_Out(add_kernel29_Valid_Out)
	);
	Batch_Norm bn_kernel29(
		.Data_A(32'b00111110110010110011111110101110),
		.Data_B(32'b00111111010000011010000001010000),
		.Data_In(add_k29_Data_Out),
		.Valid_In(add_kernel29_Valid_Out),
		.Data_Out(bn29_Data_Out),
		.Valid_Out(bn29_Valid_Out)
	);
	Relu_Core rl_kernel29(
		.Data_In(bn29_Data_Out),
		.Valid_In(bn29_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(rl29_Valid_Out)
	);
//////////KERNEL30//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111111001011001010001011010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110000001111101110100111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111101110100100001001101111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111101101011101001001110010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111101100010110000100000010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111100001100010001010101010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111110101011000010110011110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111100111101000110111000101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111101101001001010011111010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111101000110001101010010000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110100001011011001010000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111110010001101011000010111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110111000000011100101110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111110110000101001001100100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110010001101011000110000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111110000101011101011011011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111110100101101001101000011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111110010111101011001001011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111111001010000001110011101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111100000001110100011011100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110001100000110100111100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111110101101111011110101100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111110010000111111111100101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111110000110010100010111101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111110100010101101100111010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111101001111011101011011101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110110111111000110111101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110100000010011110001101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111110111110100110001110111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111101111011000101101010001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111110100001111100110011010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110100101000101110000101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111110111010110101101101001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111101111010001111011110100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111110100011011011100000010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b10111111011100111000101100101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111110100111011100101011000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111111010111001110111000100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b00111111000100111101000001010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b00111110111010110000001111011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b10111101101110100000110110010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111101110001101010001111010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111110011110010000000100111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111101001101011101101110011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111110001011001110010110100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111111000110011101100101110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b10111110101001010111111111010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111110010100100010010101111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b00111110110011001010010010100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111110011110000111000000000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b10111110001100110001110111010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111111000100001001000001100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b00111111001010011110111111010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111111100001111001010100111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b10111110100001011100111010110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b00111101000010110110000000010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b10111110011011111111001011110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b10111110001111101110000111101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111111000010011001111100111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b00111110100001001010011010101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111110100100000110011000110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b10111101001001100101001011101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111110110000011001110100101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b10111110010011000011001001011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel30_Valid_Out)
	);
	Adder_64input add_k30(
		.Data1(Data_Out_Kernel30[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel30[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel30[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel30[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel30[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel30[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel30[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel30[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel30[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel30[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel30[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel30[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel30[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel30[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel30[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel30[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel30[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel30[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel30[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel30[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel30[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel30[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel30[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel30[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel30[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel30[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel30[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel30[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel30[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel30[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel30[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel30[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel30[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel30[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel30[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel30[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel30[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel30[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel30[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel30[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel30[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel30[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel30[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel30[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel30[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel30[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel30[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel30[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel30[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel30[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel30[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel30[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel30[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel30[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel30[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel30[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel30[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel30[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel30[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel30[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel30[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel30[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel30[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel30[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel30),
		.Data_Out(add_k30_Data_Out),
		.Valid_Out(add_kernel30_Valid_Out)
	);
	Batch_Norm bn_kernel30(
		.Data_A(32'b00111110111101010101000110000001),
		.Data_B(32'b00111110110100101110110000001101),
		.Data_In(add_k30_Data_Out),
		.Valid_In(add_kernel30_Valid_Out),
		.Data_Out(bn30_Data_Out),
		.Valid_Out(bn30_Valid_Out)
	);
	Relu_Core rl_kernel30(
		.Data_In(bn30_Data_Out),
		.Valid_In(bn30_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(rl30_Valid_Out)
	);
//////////KERNEL31//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110100111110101100010000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110110011000100001000000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110010001011110110001101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110010110001110010001110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111101011011011010111000010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110110000100011000111011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111110111010111110100111101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111111001101001111000000000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111111000110000010000111010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110001101011110000011010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110110001010110110101111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111110111111010101101101011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111110100001000101010001111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111110011110011101110100101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110001101100100110111110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111101111100111011011100010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110100111000100100011001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111101000000010100111000011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110001110001100000100100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111110011001100111101101111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111111000100001100011111001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111101000100001110110111001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110101011101111001001111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111101110100010100110100110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111110001110101111001001111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111101001010100010010101110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111101110010010001001110001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110010000011000110010110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111111000011111101110010000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111110010010101000101011000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111111000110000100111011011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111110101111111111100000110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111111000000011011011100110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b00111011100011100001000110101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111111001000000000111010000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111110001001001111000110011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b10111110000011111011000100110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b00111111000010110001001010110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111110110110011001100111001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b00111111001011010110010010111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111110111011000001111001000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b10111101101011111110100001101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b00111111000100010100101011110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111100101010011101001011100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111110010011110010001101110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b10111110011110110001001000000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111110101001101101101110110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111101100101001010101010000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111111000101000010111011101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111110001011010000111110000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b10111110001111110011110101110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111110010010100101110101010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111110000110000001000001100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111110110001100100000010011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111101111010010111101111100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b00111110100010000100001110111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b10111110000000101111101000100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111110110011111110100110001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111101100010001010111011101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111111000110101010101111010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111111011110111000010001000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111110011110110110110110100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111101110010101111001101010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111110110100111010011011111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel31_Valid_Out)
	);
	Adder_64input add_k31(
		.Data1(Data_Out_Kernel31[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel31[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel31[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel31[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel31[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel31[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel31[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel31[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel31[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel31[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel31[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel31[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel31[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel31[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel31[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel31[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel31[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel31[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel31[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel31[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel31[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel31[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel31[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel31[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel31[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel31[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel31[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel31[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel31[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel31[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel31[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel31[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel31[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel31[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel31[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel31[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel31[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel31[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel31[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel31[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel31[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel31[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel31[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel31[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel31[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel31[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel31[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel31[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel31[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel31[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel31[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel31[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel31[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel31[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel31[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel31[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel31[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel31[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel31[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel31[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel31[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel31[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel31[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel31[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel31),
		.Data_Out(add_k31_Data_Out),
		.Valid_Out(add_kernel31_Valid_Out)
	);
	Batch_Norm bn_kernel31(
		.Data_A(32'b00111110111101001100000101110100),
		.Data_B(32'b10111110101010100100001101101001),
		.Data_In(add_k31_Data_Out),
		.Valid_In(add_kernel31_Valid_Out),
		.Data_Out(bn31_Data_Out),
		.Valid_Out(bn31_Valid_Out)
	);
	Relu_Core rl_kernel31(
		.Data_In(bn31_Data_Out),
		.Valid_In(bn31_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(rl31_Valid_Out)
	);
//////////KERNEL32//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111100100011111110011001111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111110000001111110010010010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110001100011101100001111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110011111101111100001110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111101011010101010011010111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111111001100000100101101000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111111000010001001111101001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111101110000100100110101000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111101101011010100000001111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111101100100001000000010000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110100000010010101010111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110100001001011001010011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110100100101001000100111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111111000010011101100111000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110011010011001101110001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111110011011101001110100010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111101000110010011111100011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111110011000000101101011001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111110101001011110001000000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111111000001011111101101011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110011101111000101110011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111111001011001110100000110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111110100100110101011011001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111101101100011101010011010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111101111100001101100000100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111101110001001011100001110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111111001010000101011010000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111101010100111011110110100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111111000100001010111001010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111101101100000011100011000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111100100100110110001111111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111110110110111100000101000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b00111110110010011111010000100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111101110110011000011001010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111110001101000110111110100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b10111110000111101111110010011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111110111100000000000100110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111110001010110110100111110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111110111010010111101111101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b00111111000000010100001001001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111111001111010101011111100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111101010110111110111010100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b00111110001001011101010110010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111111011101011110101111110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b00111110110111001001101100001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111110011010100000010110110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111111000110111111100110101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111110100000111101011111100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b00111110010101000011000111110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b00111110111101000101011101001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111101110001010100110010100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111110110001000101111011100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111101000110101000111000001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111110010011111111111010110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111111000111001010111011011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111111010000000011101010110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111111000010100110111011011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111110101011111100000110010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b10111110001110011101010111100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b00111110100110100000101101001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111101111010100110001111101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b10111110100111110010111011001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111110101110111000100101100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111110110010001001011110100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel32_Valid_Out)
	);
	Adder_64input add_k32(
		.Data1(Data_Out_Kernel32[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel32[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel32[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel32[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel32[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel32[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel32[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel32[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel32[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel32[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel32[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel32[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel32[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel32[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel32[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel32[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel32[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel32[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel32[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel32[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel32[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel32[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel32[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel32[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel32[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel32[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel32[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel32[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel32[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel32[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel32[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel32[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel32[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel32[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel32[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel32[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel32[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel32[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel32[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel32[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel32[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel32[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel32[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel32[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel32[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel32[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel32[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel32[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel32[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel32[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel32[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel32[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel32[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel32[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel32[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel32[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel32[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel32[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel32[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel32[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel32[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel32[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel32[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel32[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel32),
		.Data_Out(add_k32_Data_Out),
		.Valid_Out(add_kernel32_Valid_Out)
	);
	Batch_Norm bn_kernel32(
		.Data_A(32'b00111110111000110010110000100000),
		.Data_B(32'b00111111011011110001110110011001),
		.Data_In(add_k32_Data_Out),
		.Valid_In(add_kernel32_Valid_Out),
		.Data_Out(bn32_Data_Out),
		.Valid_Out(bn32_Valid_Out)
	);
	Relu_Core rl_kernel32(
		.Data_In(bn32_Data_Out),
		.Valid_In(bn32_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(rl32_Valid_Out)
	);
//////////KERNEL33//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111111001011011011011111100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111100101010101000110011111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110101010111100001110110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111111000111000110100001101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111110110000101001100001101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110111101111110111011001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111111011011111010101101001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111110000011111101001110000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111101101001011011100011011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111111000001010001110100101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111101100111111001111111100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110101101111000100100010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110111001110000010001011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111110101000110000110111110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110001110010011010010100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111101101010000001010001000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111011000000000000011000011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110000101010011011010110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111101010101011001000101100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111100101110010000011110001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110000011100111000001000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111101010010111010110111111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111110100111011001111011101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111101010001011001111100001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111111011101000000101111101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111110001001000010110001011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110010111011101010010110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111101110000000110100100101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111101101101100100011100000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111110110001011111000000000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111110011011000111110001101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111110100110100010100000110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111110100110011100100110100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111111000001011100011011011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111110100000000001101111010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b10111100000010111001010010001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111110010011011010010111110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111110011000110111011000001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b00111110011111110001011101101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111110110100110100110101110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111111100100001010101101110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111111000010101010011101100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b00111101010000101110110111110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b00111110001101011111101010111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b00111110111010001100110111111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b10111101101101111011111001110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111101111110000101111011111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111110110100101001111101001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111110010001110000111000110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b00111101111110101100010011000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b10111101110110000101011111010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111111000110010100011010000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111110111000100001000010001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b00111011011100110100101001000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111110111111111000101010110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b00111110100110011000011110110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b10111101010111101001101101011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111110111001101011111100100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b10111110011110001010111111010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111110101001011001001001011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111110111011010000011111101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111110101110101000011001011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b10111111000110011111011011010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b10111101101011100000001010111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel33_Valid_Out)
	);
	Adder_64input add_k33(
		.Data1(Data_Out_Kernel33[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel33[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel33[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel33[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel33[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel33[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel33[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel33[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel33[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel33[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel33[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel33[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel33[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel33[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel33[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel33[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel33[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel33[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel33[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel33[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel33[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel33[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel33[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel33[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel33[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel33[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel33[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel33[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel33[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel33[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel33[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel33[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel33[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel33[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel33[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel33[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel33[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel33[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel33[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel33[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel33[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel33[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel33[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel33[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel33[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel33[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel33[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel33[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel33[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel33[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel33[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel33[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel33[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel33[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel33[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel33[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel33[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel33[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel33[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel33[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel33[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel33[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel33[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel33[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel33),
		.Data_Out(add_k33_Data_Out),
		.Valid_Out(add_kernel33_Valid_Out)
	);
	Batch_Norm bn_kernel33(
		.Data_A(32'b00111110101111111000111011001000),
		.Data_B(32'b00111110111000000110100001011110),
		.Data_In(add_k33_Data_Out),
		.Valid_In(add_kernel33_Valid_Out),
		.Data_Out(bn33_Data_Out),
		.Valid_Out(bn33_Valid_Out)
	);
	Relu_Core rl_kernel33(
		.Data_In(bn33_Data_Out),
		.Valid_In(bn33_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(rl33_Valid_Out)
	);
//////////KERNEL34//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111101110110101110010101111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111101101101100110010101100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110110101110110111000110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110101001100110010000001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111110110110001010010111101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111110111001100110101110101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111101111110100001010111110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111010111000111011110101110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111110110001001101001101101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111110000101110101110011011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111110111010011011000100000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111110111101111000000111001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110100110000111011111001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111101111000100111100101011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110000100001010001011110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111101101110110101100010010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111111011001111111100011100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111110010011111011010011010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110001011011000111000110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111110011111010011101100011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111101101000110111011010000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111110011010001100101110111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111101110111110000000100011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111110010100111001011000010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111110111001110001001010011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111111001000111100001001011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110010110101100111100111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111101011000101101110011011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111110110010101000101100110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111110010100001111101101000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111110111000101001111011100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110100110000001100011000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111110110100111110111100000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111110110110110000011110000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111110100001110000001111110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b10111110001001010001111111101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111101000001000001101011101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111111000111001001101111101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b00111110011101111000010100100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111110000111010001010110010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b10111101001101100110101100110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b10111111000101111110001011100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111110100011001001010011010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111111000011001100010010001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b00111110110000001000111111000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111101100111010010011111111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111110010110101011000001011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111111000100100101011011011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b00111111000001101011011110001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111110110001010101100101111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111111000000001010001010010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b10111110010111110000010000010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111110000011100010000100000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111110100000011001110001001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b10111111000001111001110011000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111110110101110010101101001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b10111110011001101000101110001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111110001111000010011000000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111100101001110110000110111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b00111111000010111000100110001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111101001101110111000101000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b10111111000100000001001001000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b10111101100111000101000001000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b10111101111001101100011000010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel34_Valid_Out)
	);
	Adder_64input add_k34(
		.Data1(Data_Out_Kernel34[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel34[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel34[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel34[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel34[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel34[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel34[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel34[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel34[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel34[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel34[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel34[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel34[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel34[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel34[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel34[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel34[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel34[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel34[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel34[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel34[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel34[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel34[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel34[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel34[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel34[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel34[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel34[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel34[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel34[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel34[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel34[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel34[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel34[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel34[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel34[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel34[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel34[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel34[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel34[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel34[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel34[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel34[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel34[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel34[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel34[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel34[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel34[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel34[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel34[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel34[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel34[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel34[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel34[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel34[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel34[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel34[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel34[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel34[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel34[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel34[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel34[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel34[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel34[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel34),
		.Data_Out(add_k34_Data_Out),
		.Valid_Out(add_kernel34_Valid_Out)
	);
	Batch_Norm bn_kernel34(
		.Data_A(32'b00111110111010111100110010100111),
		.Data_B(32'b00111100110110100011100111101101),
		.Data_In(add_k34_Data_Out),
		.Valid_In(add_kernel34_Valid_Out),
		.Data_Out(bn34_Data_Out),
		.Valid_Out(bn34_Valid_Out)
	);
	Relu_Core rl_kernel34(
		.Data_In(bn34_Data_Out),
		.Valid_In(bn34_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(rl34_Valid_Out)
	);
//////////KERNEL35//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110011100100011111000000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111111000001011010011000100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110000010010001110010110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110001011010011101011100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111101001011101000001000011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111110000010100111110001110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111101101111100111001100111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111111100000010110000101010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110011010001011000110111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111110110111100010001110010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111101110011010000010101101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111101100100000101110100001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111101001000010011111101111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111110100001111100001101100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110001100101111100101101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111110011110010000011001011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111101111100001111110000110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111111000010100000111100001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110101011110100001100111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111111100000111010100100000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111111001110111010101011010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111111000000100011110011101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111110010101011100011000010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111101001000001101110101100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111110101101110011010000011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110011001101100011011101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111110011000111000010000010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111110111010010010110110101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111110001000111100110111001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111101111100001011100101100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111101110101101010100010010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111110111100010100001000101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b00111110101011101100011000111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b00111101101100011101000110110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111110101101010110110110100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b10111110010000100101110110011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111011101111010000110110101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b00111110100000010101101110001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111110000011000100011110101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111100101110011001001111010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b10111101101010011000011011000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b10111110101101101111001010000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b00111110100010011111011001001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b00111101011010111100110001111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b00111101111011111110000100101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b10111110011010101100111000010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b10111101111110110100010000110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111111100000111110000110000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b00111110001011101110100100000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111111010100110000101010101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b10111101010111000010101001010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111110000110001001011100011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b00111111000001010001010110010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111101110000110111101001111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111101011011001100011111111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111110011011010111110010000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b10111110010101110110100010000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b10111101010001111101000101001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111110110111100111111011000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111110010011101100101001011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b10111110000001110000001000000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b10111111010010110100001111011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b10111111000111111000001011000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b10111110011010010100100011010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel35_Valid_Out)
	);
	Adder_64input add_k35(
		.Data1(Data_Out_Kernel35[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel35[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel35[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel35[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel35[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel35[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel35[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel35[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel35[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel35[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel35[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel35[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel35[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel35[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel35[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel35[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel35[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel35[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel35[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel35[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel35[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel35[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel35[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel35[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel35[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel35[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel35[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel35[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel35[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel35[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel35[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel35[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel35[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel35[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel35[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel35[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel35[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel35[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel35[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel35[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel35[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel35[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel35[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel35[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel35[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel35[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel35[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel35[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel35[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel35[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel35[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel35[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel35[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel35[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel35[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel35[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel35[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel35[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel35[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel35[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel35[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel35[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel35[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel35[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel35),
		.Data_Out(add_k35_Data_Out),
		.Valid_Out(add_kernel35_Valid_Out)
	);
	Batch_Norm bn_kernel35(
		.Data_A(32'b00111110111111101000111011001111),
		.Data_B(32'b00111110111011110000111010101111),
		.Data_In(add_k35_Data_Out),
		.Valid_In(add_kernel35_Valid_Out),
		.Data_Out(bn35_Data_Out),
		.Valid_Out(bn35_Valid_Out)
	);
	Relu_Core rl_kernel35(
		.Data_In(bn35_Data_Out),
		.Valid_In(bn35_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(rl35_Valid_Out)
	);
//////////KERNEL36//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111110001011010100100010010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111100001100000000111111111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110000111000010010011011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110110011101000110111110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111110000000111001110110100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111111000001110111101111101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111110101010000110001000011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111110000001111001011111010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111110110010101111100111110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110101111100110001010100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111110110101100000000001111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110100101011001001000110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111101100001000001011010000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111110001011111010011010000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111101000001110111111001100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111110110011010100001001111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111111000111101000001100100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111011101010111010100101111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111101110000001010011110100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110111100011101011010101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111111001011111011010011000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111011111101011010000100001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110010101001100110001101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111101010010000000110011011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111101101111010011011010100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110010111000101100110111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111110001100100110011100111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110111111111001001111011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111110100000100010010011110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110101110000100111011111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111110111011110011110110111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111111000101101011010101110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b00111110110110000000110001000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111111000011111001111101100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111100000100111101010000001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111110111000000110111101011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111110011010010001000000110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b00111110000010111101100100111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111101110010000111100111111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111110100010011111000110100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111111000100111011111011111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b10111110010101101001001010110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111110001010010101000101001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111110010001100110000110110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111111000111100110111100110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b10111110000110100111111010101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111101001001010001011011010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111110111000111100001100110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111111000010001000100011000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111110110100101100101001001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111101101010010110011100010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111110000101000010011001111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111101010110011110001111000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111111000110111000100110010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111101000010011100010100000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111101110111110110010001100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b10111110100101011101001110110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b10111111001011110101101001011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b10111101111111010100101101110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b00111101001110000110011100000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b10111110001001010000011000011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111110100010011010110010101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b10111111100110111010100110100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b10111111000100111101010000110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel36_Valid_Out)
	);
	Adder_64input add_k36(
		.Data1(Data_Out_Kernel36[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel36[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel36[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel36[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel36[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel36[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel36[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel36[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel36[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel36[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel36[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel36[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel36[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel36[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel36[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel36[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel36[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel36[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel36[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel36[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel36[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel36[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel36[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel36[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel36[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel36[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel36[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel36[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel36[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel36[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel36[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel36[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel36[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel36[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel36[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel36[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel36[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel36[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel36[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel36[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel36[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel36[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel36[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel36[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel36[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel36[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel36[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel36[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel36[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel36[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel36[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel36[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel36[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel36[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel36[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel36[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel36[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel36[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel36[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel36[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel36[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel36[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel36[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel36[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel36),
		.Data_Out(add_k36_Data_Out),
		.Valid_Out(add_kernel36_Valid_Out)
	);
	Batch_Norm bn_kernel36(
		.Data_A(32'b00111110111110100010100100100010),
		.Data_B(32'b00111111010010011001001111010101),
		.Data_In(add_k36_Data_Out),
		.Valid_In(add_kernel36_Valid_Out),
		.Data_Out(bn36_Data_Out),
		.Valid_Out(bn36_Valid_Out)
	);
	Relu_Core rl_kernel36(
		.Data_In(bn36_Data_Out),
		.Valid_In(bn36_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(rl36_Valid_Out)
	);
//////////KERNEL37//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110011101000001001001001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110001000101001001000001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110100101100100001110010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111101101101101010110010000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111101110110010011001000011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111100001001000011110101101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111111001111100100010001100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111110001001101101010001110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111101011100101111001110001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111101010001001100000001110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111100101100111110110001101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110001100101101111011110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111110101100101011100111101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111101111111100000001010001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111111000010011001100101111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111110011001110001100010101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111110011110000010000110010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110101010011001010101100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111101100001000111100101100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111110110111111000010010110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111111001110110010010110010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111101010000101110100100110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110010110100000100111010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111110011100110101110011100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111110101000000000001111010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110011000001111111011001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111101111101111010101001111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111110100100100000010111001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111110101010000001010011010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110011010110000011011111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111111000010100101010111111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111111011110111000000111001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b00111111001011010111111011000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b00111110000010010100000111000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111101111000100011111011001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b10111100001110101010101010010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b10111110100011010100001101010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111100000111000100111011000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111111001110111110010001001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111110111001110000010100011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111110110111000001000011001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b10111110110001111100010101011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b00111110010011101100111010010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111110001000110111101000000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b00111110000011001000101001100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111111001001101010001000001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b10111110010001010110101010111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b00111100000010101110010011011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111101001101001110010111111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b00111111010001000110001100100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111110111001100101111100010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b10111111000100101110000100011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b00111110000101000000000101001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111111000000110011011110110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111110000110010000001101011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111110111001011101001011111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b10111101110000111001110011000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111110100110011011100011001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111110010100000101001100111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b00111110011001101111110111010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111111000010110110100000110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111110101100110011101110010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111110101001110001110010111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b10111110111001000000110100000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel37_Valid_Out)
	);
	Adder_64input add_k37(
		.Data1(Data_Out_Kernel37[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel37[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel37[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel37[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel37[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel37[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel37[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel37[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel37[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel37[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel37[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel37[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel37[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel37[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel37[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel37[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel37[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel37[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel37[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel37[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel37[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel37[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel37[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel37[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel37[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel37[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel37[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel37[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel37[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel37[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel37[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel37[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel37[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel37[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel37[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel37[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel37[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel37[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel37[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel37[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel37[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel37[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel37[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel37[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel37[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel37[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel37[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel37[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel37[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel37[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel37[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel37[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel37[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel37[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel37[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel37[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel37[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel37[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel37[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel37[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel37[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel37[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel37[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel37[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel37),
		.Data_Out(add_k37_Data_Out),
		.Valid_Out(add_kernel37_Valid_Out)
	);
	Batch_Norm bn_kernel37(
		.Data_A(32'b00111111000001100011010110000001),
		.Data_B(32'b00111110111010001101111000010000),
		.Data_In(add_k37_Data_Out),
		.Valid_In(add_kernel37_Valid_Out),
		.Data_Out(bn37_Data_Out),
		.Valid_Out(bn37_Valid_Out)
	);
	Relu_Core rl_kernel37(
		.Data_In(bn37_Data_Out),
		.Valid_In(bn37_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(rl37_Valid_Out)
	);
//////////KERNEL38//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111111000001110001111111100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111110000010100001110001010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111101011110110110000000001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110010010101110101000100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111110101011010011000011001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111110001001001001010110001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111110110110010101101001000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111110100110101000110011100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110100110001001010000100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110101101110111100111110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110000010001100100100010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111111000000111000001010001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110100101010110100101011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111110001111000011100001110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111101111010101111101010101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111110011100110111011101101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111110100001001111010100011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111100101100110000111110110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110001110110100101101010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110111001000011010000011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110000010100011100110001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111111001000110101110100111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111111010100111001000010000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111101100101011111111111011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111110000010000111110100011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111100010000011100110011100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110000101011001100110100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110011110110110010011110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111100101001010110000101101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111110001100110010001010101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111101101101011110010100001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111101000011000000011110010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b00111110110011010001011101111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111110101011010111010100001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111100001111110110001011011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111111101000010000110011011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b10111101010001101001111100101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b00111101010111001000011100100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b00111110101111010010010010010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b00111110010000001100111110111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111110010011000101000011101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b10111101110100010000000111011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b00111110000000011010111101101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b00111110100100110010010101100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b00111101111010110111011110001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111110011100010101110000111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b10111110111100011100111111111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111111001011001000000000000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b00111111010000111010001001111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b00111110010101101100100110100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111110110000110111011011110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b10111111000100000101110111011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b00111110110010000010111000100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b00111101000000100000110100001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111110100101101110001111001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111110100000001110000010011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b10111110111100001111000101110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111101101010101011001111011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b10111110000001100101101011110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111111000100001101101100111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111110101111100010000111111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111100011001000011110011110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111001111111110000101000001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b10111101110000101101001110000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel38_Valid_Out)
	);
	Adder_64input add_k38(
		.Data1(Data_Out_Kernel38[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel38[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel38[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel38[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel38[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel38[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel38[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel38[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel38[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel38[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel38[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel38[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel38[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel38[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel38[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel38[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel38[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel38[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel38[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel38[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel38[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel38[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel38[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel38[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel38[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel38[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel38[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel38[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel38[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel38[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel38[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel38[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel38[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel38[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel38[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel38[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel38[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel38[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel38[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel38[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel38[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel38[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel38[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel38[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel38[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel38[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel38[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel38[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel38[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel38[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel38[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel38[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel38[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel38[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel38[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel38[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel38[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel38[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel38[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel38[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel38[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel38[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel38[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel38[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel38),
		.Data_Out(add_k38_Data_Out),
		.Valid_Out(add_kernel38_Valid_Out)
	);
	Batch_Norm bn_kernel38(
		.Data_A(32'b00111110111001001001100000100100),
		.Data_B(32'b00111111000001101010110111010000),
		.Data_In(add_k38_Data_Out),
		.Valid_In(add_kernel38_Valid_Out),
		.Data_Out(bn38_Data_Out),
		.Valid_Out(bn38_Valid_Out)
	);
	Relu_Core rl_kernel38(
		.Data_In(bn38_Data_Out),
		.Valid_In(bn38_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(rl38_Valid_Out)
	);
//////////KERNEL39//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111110000011100000011100010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110101110111110100001100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111101011000100000101001000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111111001001100011111011011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111101000000101011011110000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111110100001011110101101110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111111100000001111110110110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111011110110001101111001111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111101110111011110011111101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110100110101101001010110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111110110110001001001001011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110100001001100011101110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111111000001000101011011011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111110100110011111000111001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111101011001111011110000111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111110101111100011010000100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110101110101101100000011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111101010011011111100010001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110111100101110100101000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111110100100110110000110101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110000111110011010111000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111101101101111101110101100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111101001110110010111100000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111110000110011011101101001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111101111111001101111001110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110110101101000100000111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111111000111110100101010000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111110001000111101110010011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111110001100000001110000101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111101001011010111100110100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111101100111000000100011011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111110101110100011010001101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b00111110011100010110001110010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b00111110010100010010011100010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111101010011100010001101011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b10111110101010110111011100111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b10111110010110010100011110000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b00111101001010110111010001000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111110101101000001110100101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111110110011011110101100101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111110110000111010101001010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b10111101011001110110111000111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111110111010011100010011110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b00111111001011010000010010100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111111000101001000010011001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111100001110110101001100101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111110001101100011101011110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b00111110101101011110100001101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b00111101011111000111101111010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b00111110100110110000111100101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b10111111000100001111100101010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111110001010111111011010011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b00111110010011000011110001011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b00111110100111111011100001100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111111001101111010101101010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111101100011001100110011010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b10111110001000110100010110101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111111001100100100101010100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b10111100100000111011101011111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111111000101110011100001100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111100010000100111010101100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b10111110111111100101101110110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b10111110101111100101001001000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b10111111000000011100001010001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel39_Valid_Out)
	);
	Adder_64input add_k39(
		.Data1(Data_Out_Kernel39[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel39[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel39[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel39[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel39[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel39[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel39[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel39[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel39[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel39[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel39[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel39[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel39[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel39[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel39[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel39[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel39[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel39[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel39[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel39[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel39[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel39[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel39[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel39[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel39[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel39[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel39[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel39[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel39[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel39[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel39[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel39[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel39[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel39[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel39[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel39[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel39[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel39[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel39[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel39[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel39[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel39[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel39[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel39[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel39[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel39[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel39[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel39[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel39[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel39[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel39[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel39[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel39[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel39[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel39[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel39[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel39[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel39[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel39[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel39[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel39[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel39[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel39[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel39[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel39),
		.Data_Out(add_k39_Data_Out),
		.Valid_Out(add_kernel39_Valid_Out)
	);
	Batch_Norm bn_kernel39(
		.Data_A(32'b00111110111111101101110000110111),
		.Data_B(32'b00111110110110111100101100001100),
		.Data_In(add_k39_Data_Out),
		.Valid_In(add_kernel39_Valid_Out),
		.Data_Out(bn39_Data_Out),
		.Valid_Out(bn39_Valid_Out)
	);
	Relu_Core rl_kernel39(
		.Data_In(bn39_Data_Out),
		.Valid_In(bn39_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(rl39_Valid_Out)
	);
//////////KERNEL40//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110010111111001011011011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111101111000000011110110110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110001111010101001101110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111101100010100011000010011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111111000110110110110101000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111100001100111110111100110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111111000001101010000010101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111110011000010110001101110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110010001001111010111001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111011101011001110011100001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111110001011100101010101111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111101100101001011000001001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110000000101010100100100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111111000111110111111100011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110111000111001011001010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111110111001101011101101100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111110111001000111110110010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110111010001111110010010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111110110101100101011100110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111110100101010001001001101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110110000001110010000110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111111011111001100010111001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111110110100000110001011111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111110100010101000010101011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111110001100101111010010100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111111000101111101011101000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111110010011101100000000000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110010100110010110110110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111110110010000111101011101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111101110110010001000110001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111110011011010111001101010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111110011000111101111011010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b00111111000010110001101111001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111110100100110010010010100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111110111010001101110010010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b10111100111110110011011010110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111111000000111100010000011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b00111110000000100110011001000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b00111110111101100011111010011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b00111110010000000010100110000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b10111110001111111101000001010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b10111110101111011100101111100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111110100101101011101010100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b00111111010010111011111000111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b00111111000101011100100110110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b10111110001011110101101110101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b10111110100001010000010000111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111111001101111100101111100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b00111110000001011001001010000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111110111100100100000000101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111110001011110000001010100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b10111110010001101000001110010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b00111101011101100111111100000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111110101111000101110010001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111110010001110010001000000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111101101001111111101101000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111110001011011011111010001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111111001011101100110110100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111101100001110001001111101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111110100010000110001110001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111110110100110101100111001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b10111101101000001010111110100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111101110001010001010111000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111111001000111101001010001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel40_Valid_Out)
	);
	Adder_64input add_k40(
		.Data1(Data_Out_Kernel40[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel40[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel40[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel40[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel40[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel40[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel40[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel40[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel40[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel40[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel40[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel40[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel40[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel40[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel40[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel40[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel40[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel40[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel40[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel40[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel40[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel40[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel40[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel40[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel40[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel40[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel40[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel40[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel40[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel40[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel40[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel40[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel40[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel40[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel40[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel40[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel40[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel40[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel40[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel40[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel40[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel40[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel40[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel40[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel40[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel40[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel40[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel40[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel40[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel40[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel40[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel40[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel40[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel40[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel40[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel40[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel40[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel40[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel40[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel40[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel40[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel40[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel40[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel40[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel40),
		.Data_Out(add_k40_Data_Out),
		.Valid_Out(add_kernel40_Valid_Out)
	);
	Batch_Norm bn_kernel40(
		.Data_A(32'b00111110111010011011101010010011),
		.Data_B(32'b00111111010011101011111010001011),
		.Data_In(add_k40_Data_Out),
		.Valid_In(add_kernel40_Valid_Out),
		.Data_Out(bn40_Data_Out),
		.Valid_Out(bn40_Valid_Out)
	);
	Relu_Core rl_kernel40(
		.Data_In(bn40_Data_Out),
		.Valid_In(bn40_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(rl40_Valid_Out)
	);
//////////KERNEL41//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110100011111111101000000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110110110111011010101111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110000100010100110111000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110110111000111001010111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111111001011101110100001101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111110101110000110111111001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111101111100000111001000011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111110101110000100001110111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111101110111110101001101001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111110111111110000111011100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110010011010010010101001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111110010000111100100101000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110011111101010011011000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111110101011000101010111100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110000001010111000111010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111110101111001100111111000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111110110100000110000100010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111110100011011011011111011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110011101010101110111110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110110101001010101101110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111100111110111001101101110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111110111000111011011111110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110100110111111110011001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111100000001101111101001111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111101111011001111100110100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110010000000001100100001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111111010010001010101001111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110110101011110010001100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111110101101011111101110101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111110001100101111111000111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111101101010010010000011110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111110000101101111011111000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b00111110001000110001100111011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111111000111110010110010000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111111000100111101110000110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111110111001101111110100000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b10111110110001111010111101001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b00111110110001001101100100000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b00111111100111101010000111000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111011010100010001111101101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111110110111011101100011000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b10111110001000011011001000010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b00111110011000100010011101011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111101110101011000111011011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111110000010101010001101101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111100101010101110111101100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111110010101011110001000100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111101010111001101111101011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111110101101010001010011110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111110000100101010011101011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b10111110100010001001011000111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b10111110100011000111001110101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111101011001010010010001001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111111001110111011011011011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111101111110011100011000000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111111001011111100110100110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111101011101110100111111111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b10111110101101000010011110101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b10111111000010000001011011010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111100100010110010100101010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111110010101100101111000110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111110000100100001000000110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111101011111000110000000011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111110000010011010101011101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel41_Valid_Out)
	);
	Adder_64input add_k41(
		.Data1(Data_Out_Kernel41[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel41[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel41[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel41[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel41[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel41[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel41[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel41[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel41[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel41[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel41[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel41[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel41[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel41[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel41[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel41[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel41[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel41[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel41[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel41[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel41[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel41[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel41[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel41[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel41[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel41[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel41[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel41[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel41[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel41[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel41[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel41[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel41[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel41[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel41[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel41[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel41[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel41[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel41[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel41[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel41[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel41[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel41[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel41[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel41[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel41[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel41[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel41[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel41[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel41[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel41[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel41[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel41[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel41[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel41[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel41[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel41[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel41[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel41[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel41[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel41[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel41[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel41[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel41[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel41),
		.Data_Out(add_k41_Data_Out),
		.Valid_Out(add_kernel41_Valid_Out)
	);
	Batch_Norm bn_kernel41(
		.Data_A(32'b00111110110101110011011111110000),
		.Data_B(32'b00111110100111110000100001110001),
		.Data_In(add_k41_Data_Out),
		.Valid_In(add_kernel41_Valid_Out),
		.Data_Out(bn41_Data_Out),
		.Valid_Out(bn41_Valid_Out)
	);
	Relu_Core rl_kernel41(
		.Data_In(bn41_Data_Out),
		.Valid_In(bn41_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(rl41_Valid_Out)
	);
//////////KERNEL42//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111101101011110000011100110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111101001011110110110000001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111111000100111101111111100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110111011011010000000100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111101111110000010010110100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111101110001010111101000101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111101101011001100001010110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111110100111000010110101101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111110110001100011010001000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110100110001100100001111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111110010100000110110000110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111100001110110010000011010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111101000000000111010000010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111111000110101110111011110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111101101011001110101001011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111111000000101001011110100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111101111101111010100111110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111110100011010101101101010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111110100111100111000010101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111111100000011001110001101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110110000001001111011110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111101111001010101010110000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111111001011011111111001010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111110001101101101010001010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111010000010101111100001000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110100010111000011110100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111101100000100111110100110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111100100010010010010000111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111110110010000001111011111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110000100101100101001011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111110101000011100111111011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110001001111010111111001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b00111101101010110110001100101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b00111110001110101001000111100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111110100111010000001101110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111111010111011000001111111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111110111110001111101011001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b00111101101011001100001001110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b00111111000101100000001000100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111110000101000010011000101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111011010010110110110010111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111110110011001000111110110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b00111110111100000001110011101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111110011110111101000000001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111111000100011010001011100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b10111111000000011011111100001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111110000011001101101100101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b00111110100101110110111010111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111111000001001010101111000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b00111110111101101111000110111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111101000101111110100011111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111101111100101000100010101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b00111101010111100110010100011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b00111111001001000110101001011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111110001011000101001001110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111110011010110000001000100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b10111110000101000011100100011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111101010101100010101100001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111101100011000101011010100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111101110110001101010011110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111111010000001110110001110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b10111110000100010100000111100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b10111111001110100000111100000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b10111111000101101100000100101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel42_Valid_Out)
	);
	Adder_64input add_k42(
		.Data1(Data_Out_Kernel42[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel42[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel42[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel42[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel42[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel42[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel42[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel42[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel42[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel42[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel42[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel42[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel42[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel42[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel42[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel42[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel42[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel42[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel42[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel42[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel42[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel42[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel42[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel42[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel42[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel42[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel42[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel42[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel42[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel42[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel42[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel42[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel42[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel42[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel42[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel42[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel42[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel42[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel42[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel42[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel42[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel42[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel42[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel42[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel42[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel42[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel42[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel42[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel42[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel42[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel42[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel42[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel42[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel42[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel42[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel42[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel42[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel42[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel42[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel42[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel42[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel42[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel42[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel42[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel42),
		.Data_Out(add_k42_Data_Out),
		.Valid_Out(add_kernel42_Valid_Out)
	);
	Batch_Norm bn_kernel42(
		.Data_A(32'b00111110111001101111111001010111),
		.Data_B(32'b00111101111111100001011001111001),
		.Data_In(add_k42_Data_Out),
		.Valid_In(add_kernel42_Valid_Out),
		.Data_Out(bn42_Data_Out),
		.Valid_Out(bn42_Valid_Out)
	);
	Relu_Core rl_kernel42(
		.Data_In(bn42_Data_Out),
		.Valid_In(bn42_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(rl42_Valid_Out)
	);
//////////KERNEL43//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111110011110100110100111110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110101000110011001110001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110101100001000110001101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110000101000010010110101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111110100001101001110111100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110001101001011011010110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111111000000110000110001000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111110111010111100011101011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110100101001101011100011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111101100110000011111000110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110010111110010000000001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111110100010010110001101010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110011110101101001100111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111110101011011010111110001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110011110111001111011100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111110011000100000111110101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111111000001001001101101111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111110010111000001010100000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111101110100100111011100000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110100101111110010100111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111111000010101101001101000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111110110011000101110001011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111101111010000110011011111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111100110110011001100110001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111110110111000101010110011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111111000001001010101000101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110010100111110010000001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111101101101010001111001100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111101110000100000110001010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111111001100110010110010101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111111000111000010111100011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111110011011101010010010000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b00111110000000001100100011010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111111000011110000111111001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111111000011001001111100010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111110011010101000100000001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111111010001100101011010111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111101101010001111011011000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b00111110000101001011100010110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b00111101110001110111101011000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b10111110101101100110110011010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111110100010010100011000011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b00111110111111100010010111101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111110011010010000100111000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111111000010110101001000011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111110100100100101000011010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b10111110010001010010000111001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b00111110010000100111110001011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b00111110111000110001000001001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b00111101111111110001101001111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b10111110100100001010100110011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111110101011110101001101100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111110100010001011011111000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b00111110111001000010100010111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b10111101100000010101011101111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b00111101000011001001110111000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111110111100001110110111111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111110001010010011001100010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b10111110001011111111000010010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b00111110000010010110110001011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111110110000111100010111110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111111001101010001000101111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b10111110010111101100010011101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b10111111010000011101110010001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel43_Valid_Out)
	);
	Adder_64input add_k43(
		.Data1(Data_Out_Kernel43[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel43[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel43[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel43[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel43[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel43[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel43[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel43[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel43[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel43[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel43[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel43[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel43[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel43[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel43[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel43[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel43[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel43[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel43[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel43[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel43[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel43[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel43[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel43[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel43[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel43[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel43[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel43[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel43[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel43[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel43[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel43[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel43[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel43[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel43[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel43[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel43[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel43[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel43[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel43[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel43[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel43[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel43[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel43[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel43[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel43[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel43[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel43[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel43[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel43[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel43[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel43[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel43[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel43[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel43[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel43[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel43[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel43[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel43[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel43[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel43[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel43[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel43[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel43[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel43),
		.Data_Out(add_k43_Data_Out),
		.Valid_Out(add_kernel43_Valid_Out)
	);
	Batch_Norm bn_kernel43(
		.Data_A(32'b00111111000010000110001000110110),
		.Data_B(32'b00111110111110110001101011000110),
		.Data_In(add_k43_Data_Out),
		.Valid_In(add_kernel43_Valid_Out),
		.Data_Out(bn43_Data_Out),
		.Valid_Out(bn43_Valid_Out)
	);
	Relu_Core rl_kernel43(
		.Data_In(bn43_Data_Out),
		.Valid_In(bn43_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(rl43_Valid_Out)
	);
//////////KERNEL44//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111101101010011101111101111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111101101110010110001110101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110000010100100101000010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110001011011000011110110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111110100010011110000011111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110010011001000110100001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111101111100111101111110111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111111000111111010101001000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110100111111111000101010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111111000110011011010010000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111101011110111111101001001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111101010001011101000100110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110010111000110100010000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111110110110011010001001011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111101000010111010000011000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111110100010111011000000100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111111001011001000111001110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111110010011101011011100011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111101110001011110011010011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111110111110110110010110001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110111011111010101001010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111110110001010011100111000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111111001100111000010001101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111110111000101100100011101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111110000110010011011001100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111101001010000011001001111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111111000111011101110001110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110110110110000000011000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111110001010000011101101000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111100111110001011011111000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111111000011010100000111000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111101010111100100110010010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111101010000001110100110011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111101111010100100101011100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111110011010001101011010101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111101100011001110110010011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b10111110110000101000111111111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b00111110011101101111001000100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111110010000001110101011100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111101111100001010011111100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b10111110100001000110111011111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b10111110111010001100101000011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b00111111001010101100000011011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111101000001010000101101001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111111100101000011011111110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b10111111010100010001111111111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b10111110010001000000100011010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b00111110110011101100111001100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b00111110110110011000100010001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b00111110100000000001100101110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b10111110111100010000110000010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b10111011111011010000111110110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111110010000001101001110001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111110110000000101111101101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111110011001111001111010000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111110110101000000111011111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b10111110101000000001000010110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b10111110100110100100000111010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111110101110101100101010101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111110110001011011111001101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b10111100110100110110110001110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b10111110101001011000110010111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111110011010010000011110111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b10111101100101011010010101000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel44_Valid_Out)
	);
	Adder_64input add_k44(
		.Data1(Data_Out_Kernel44[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel44[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel44[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel44[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel44[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel44[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel44[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel44[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel44[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel44[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel44[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel44[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel44[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel44[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel44[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel44[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel44[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel44[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel44[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel44[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel44[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel44[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel44[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel44[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel44[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel44[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel44[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel44[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel44[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel44[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel44[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel44[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel44[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel44[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel44[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel44[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel44[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel44[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel44[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel44[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel44[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel44[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel44[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel44[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel44[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel44[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel44[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel44[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel44[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel44[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel44[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel44[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel44[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel44[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel44[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel44[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel44[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel44[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel44[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel44[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel44[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel44[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel44[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel44[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel44),
		.Data_Out(add_k44_Data_Out),
		.Valid_Out(add_kernel44_Valid_Out)
	);
	Batch_Norm bn_kernel44(
		.Data_A(32'b00111110110111101010000111011000),
		.Data_B(32'b10111100101001100000011110100001),
		.Data_In(add_k44_Data_Out),
		.Valid_In(add_kernel44_Valid_Out),
		.Data_Out(bn44_Data_Out),
		.Valid_Out(bn44_Valid_Out)
	);
	Relu_Core rl_kernel44(
		.Data_In(bn44_Data_Out),
		.Valid_In(bn44_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(rl44_Valid_Out)
	);
//////////KERNEL45//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111101110011111110000101001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111111000010100000010001100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111101001100010010100000101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110100001010110110100101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111110010011100010100111001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110001100110111000100000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111111011000010101011001110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111110110100110011100110101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110100100101100001101011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110100111001010101011011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111101001010011100010101110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111111010100001111001110010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111011011010100010100000111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111111001111001100110000100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111111010000110010011111111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111101001000110000001110001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110101100011011010111110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111101001010111010100110010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110001101011100010000001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111101101110101000111011010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111111000000011111111011011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111111011000000110000111111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110100101000111010111110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111110100101001001011001110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111110000100100111110101111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111101100001001111001011100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111110100001110110110110000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111101101000011111110101010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111101111001110001101001001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111111001010100111100111110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111110100100010111101011100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111100000110000100001000011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111110101100011110000100110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111110000101010111000101110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111101110000111111100110001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111110111110111100100110111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111111001010010000010001011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b00111111000010000111100000011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b00111101000110101110011010101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111110100100001011100000001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111101110110111101111110100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b10111110110000110000110001000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111110110101011101110111110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111101100100100001010100000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111110010001001010110001101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b10111111001001111010011000110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b10111110100001010110100111110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b00111101011111101110101010101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b00111110000100000100111001000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b00111110010110000110101111000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111010100011010101001000001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111111001001110110010101001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111110011111011010101101001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111111000110110101101010110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111111000000011000001101000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111100010111001001101111000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111110100010010010100100001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111100110100101010100000000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b10111101010011101001110110111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b00111110110101100011100010110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b10111100010101000001110000010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b10111100011010010010110011101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111110110010101010110011110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111101100011111110001111111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel45_Valid_Out)
	);
	Adder_64input add_k45(
		.Data1(Data_Out_Kernel45[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel45[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel45[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel45[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel45[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel45[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel45[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel45[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel45[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel45[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel45[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel45[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel45[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel45[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel45[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel45[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel45[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel45[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel45[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel45[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel45[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel45[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel45[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel45[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel45[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel45[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel45[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel45[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel45[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel45[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel45[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel45[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel45[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel45[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel45[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel45[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel45[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel45[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel45[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel45[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel45[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel45[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel45[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel45[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel45[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel45[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel45[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel45[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel45[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel45[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel45[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel45[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel45[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel45[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel45[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel45[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel45[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel45[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel45[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel45[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel45[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel45[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel45[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel45[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel45),
		.Data_Out(add_k45_Data_Out),
		.Valid_Out(add_kernel45_Valid_Out)
	);
	Batch_Norm bn_kernel45(
		.Data_A(32'b00111110111001000010000110010100),
		.Data_B(32'b00111111000101010110011110110111),
		.Data_In(add_k45_Data_Out),
		.Valid_In(add_kernel45_Valid_Out),
		.Data_Out(bn45_Data_Out),
		.Valid_Out(bn45_Valid_Out)
	);
	Relu_Core rl_kernel45(
		.Data_In(bn45_Data_Out),
		.Valid_In(bn45_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(rl45_Valid_Out)
	);
//////////KERNEL46//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111101000000111010110110000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111101100111111110100111101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111101101101000010001010110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110010000110101010101100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111110100100000100110110111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111101100001100001111110010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111110100101001101001110110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111101011110010010001110111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111101111001101000001101101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111110011110011110011111010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111101010000111110111010010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111101100010111100011111101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111101111011001010000000111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111011110010100111101110100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110010000111100010111110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111110000100111010011010111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111101000010101001001110000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110010111000111111011101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111111100011010010100010110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111111011101100101001000111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110101001101110000010000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111101100111111100101011010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110001011000101101001100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111110001111001110011111011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111011101100010000101010010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110011110011111010100000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111110000100001010100011010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111101011100100101001001100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111101110100100111010001101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111111000100110001010111100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111110110011010011001001001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111110000111111010110111000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b00111111000100100001000101010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111111001111010110000010010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111110001000011000101101010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b10111101010000110010100101011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b10111111001000110101010100010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111110110000110100111101010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b00111111000010000010000110000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b00111110101111011101011000100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111110010111111010010010010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b10111101100000101100111000100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b00111101000100001001011100100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b00111110011111000101101110110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111110101111101010010010111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b10111101011110000001000100000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111110001001001111011101111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111111001000110100101100111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111101010001011111011011101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111111001001111000000011010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b10111110000101101000000100111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111111011100000100100101001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b00111111001100111011010101011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b00111110101000010010110011000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111110110100001110111100001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111110111000001011010111000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b10111110100010011011011110011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111110101100011000110010101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111110111000010000101011011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111110101110001111101110110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111101000101100110110011111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b10111110111100100100110011110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111110100001011001111111101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111110100101011010000011110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel46_Valid_Out)
	);
	Adder_64input add_k46(
		.Data1(Data_Out_Kernel46[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel46[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel46[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel46[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel46[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel46[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel46[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel46[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel46[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel46[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel46[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel46[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel46[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel46[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel46[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel46[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel46[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel46[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel46[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel46[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel46[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel46[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel46[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel46[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel46[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel46[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel46[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel46[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel46[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel46[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel46[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel46[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel46[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel46[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel46[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel46[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel46[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel46[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel46[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel46[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel46[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel46[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel46[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel46[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel46[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel46[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel46[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel46[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel46[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel46[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel46[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel46[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel46[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel46[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel46[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel46[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel46[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel46[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel46[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel46[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel46[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel46[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel46[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel46[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel46),
		.Data_Out(add_k46_Data_Out),
		.Valid_Out(add_kernel46_Valid_Out)
	);
	Batch_Norm bn_kernel46(
		.Data_A(32'b00111110110100000110100010001101),
		.Data_B(32'b00111111001000011110101101100100),
		.Data_In(add_k46_Data_Out),
		.Valid_In(add_kernel46_Valid_Out),
		.Data_Out(bn46_Data_Out),
		.Valid_Out(bn46_Valid_Out)
	);
	Relu_Core rl_kernel46(
		.Data_In(bn46_Data_Out),
		.Valid_In(bn46_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(rl46_Valid_Out)
	);
//////////KERNEL47//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111101010000101000100101100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111110100001011101011110101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110110010011000111101001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110001010010010000001101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111110111000110011111110000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111111000011100100101011010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00110111110000010100001111010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111111001110000010000100110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110100110101100110100100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110110100101100011011000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111110001100010011000000101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110011100000010010000100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111110011101011111111010010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111110100110000011001000101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111111001110000111000101100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111111000001011011111100100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110100000000111011110101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110100001101010000011000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111111001000110000111010011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111100010010100000011001011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110000111010001011100100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111111000101101100110110111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111110010101011101100000111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111111000011000100110101000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111111010110001100101110010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110101011010001100010001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110001010011011010110100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111101100001101010110000001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111111000001011100001100111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110101110011101011111000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111101101100011111011111111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111101000011010011001001001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b00111101010011000011001110001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b00111110000101101110011001000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111110011101011001010001111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111110101100100000100001011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111110001101001111110010010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111110010100001100100101000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b00111110100001010001011100000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111101011100010010011011010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b10111111000011111011110011100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b10111111001101101100010001000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b00111110101111000101010100110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b00111110101000111011000000011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111111000000011000101011111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111111010000100110111011001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b10111110100000100010111000110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b00111110111000100111010001010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111101100110111000110110001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111100001000111000101000010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b10111110010001011001101101010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111111000100000101111001011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111100100111000110101001100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111101100111001011110000011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b10111101100010001110110110101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111101000100011010100000100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b10111101101100100110101001010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b10111110100000111100001010101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b10111110110011001100011101011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b00111101111101011111001001101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111101000110111001010111111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111110001100110100101000010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111110111010010111001111001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111111010010101100010111001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel47_Valid_Out)
	);
	Adder_64input add_k47(
		.Data1(Data_Out_Kernel47[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel47[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel47[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel47[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel47[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel47[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel47[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel47[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel47[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel47[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel47[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel47[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel47[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel47[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel47[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel47[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel47[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel47[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel47[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel47[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel47[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel47[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel47[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel47[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel47[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel47[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel47[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel47[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel47[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel47[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel47[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel47[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel47[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel47[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel47[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel47[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel47[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel47[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel47[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel47[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel47[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel47[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel47[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel47[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel47[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel47[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel47[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel47[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel47[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel47[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel47[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel47[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel47[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel47[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel47[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel47[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel47[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel47[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel47[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel47[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel47[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel47[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel47[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel47[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel47),
		.Data_Out(add_k47_Data_Out),
		.Valid_Out(add_kernel47_Valid_Out)
	);
	Batch_Norm bn_kernel47(
		.Data_A(32'b00111110110110000001000100100100),
		.Data_B(32'b00111110101111111110000000011011),
		.Data_In(add_k47_Data_Out),
		.Valid_In(add_kernel47_Valid_Out),
		.Data_Out(bn47_Data_Out),
		.Valid_Out(bn47_Valid_Out)
	);
	Relu_Core rl_kernel47(
		.Data_In(bn47_Data_Out),
		.Valid_In(bn47_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(rl47_Valid_Out)
	);
//////////KERNEL48//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110001101110100110011100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111111001100111010001110100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110001110111101010111000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111101111001100111101100011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111101101111011101001011011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111110101111101011111011110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111101101011100111110001110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111110100011000111111111101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111101000001010111100011000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111110000111010000100010001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111110101000001000101100010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111101100110111000001001101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111111001010111001110001001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111101110011011010001111011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110100001111110001011001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111101011100100000000011011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110100011100000011101010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111110101001000011111100111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111111000011100000000100111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111101100100010000110100010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111100110001011111110010000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111110111010100001101111111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111110001110000100001001000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111101001110101001000101011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111111000101111101100111111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111101100010001100101110101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111101100011110100010011101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110000110110010111011000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111110011001000010011011001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111100000100001000010011101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111111011010010101111100101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110011000000010101001100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111110100000100111011011000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b00111100100101010110000100001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111101110100100001000010010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b10111110100010111011111001000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111101111011010111000000101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111110100100100000001110110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111110101010001110011010000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111110111100010010110111001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111110000010011100010110110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111111001100011011010100111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111111000001100010110110111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111110101010000010110010011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b00111110010100010110000001101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111100010111110010011101011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111111001000000101111110101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b00111101110111000100111001100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b00111111000011000100001111001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111110100110101001101000010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b10111110110101011101111100001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111101111000010010111100100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111100110101111101000101101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111101110001000011101110001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111110110000111100111111000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111110111001110111001001111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111111001000111001101011100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111101011011011100010001110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111101100101000000110001110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b00111111001000101110101000001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111110000010101100000100101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111111001100110110110100100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111111010110001001101001011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111110110100000011100010000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel48_Valid_Out)
	);
	Adder_64input add_k48(
		.Data1(Data_Out_Kernel48[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel48[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel48[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel48[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel48[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel48[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel48[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel48[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel48[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel48[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel48[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel48[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel48[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel48[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel48[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel48[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel48[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel48[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel48[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel48[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel48[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel48[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel48[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel48[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel48[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel48[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel48[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel48[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel48[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel48[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel48[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel48[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel48[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel48[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel48[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel48[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel48[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel48[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel48[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel48[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel48[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel48[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel48[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel48[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel48[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel48[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel48[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel48[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel48[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel48[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel48[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel48[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel48[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel48[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel48[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel48[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel48[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel48[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel48[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel48[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel48[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel48[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel48[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel48[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel48),
		.Data_Out(add_k48_Data_Out),
		.Valid_Out(add_kernel48_Valid_Out)
	);
	Batch_Norm bn_kernel48(
		.Data_A(32'b00111110110111001101001001000100),
		.Data_B(32'b00111111001000011100110100101010),
		.Data_In(add_k48_Data_Out),
		.Valid_In(add_kernel48_Valid_Out),
		.Data_Out(bn48_Data_Out),
		.Valid_Out(bn48_Valid_Out)
	);
	Relu_Core rl_kernel48(
		.Data_In(bn48_Data_Out),
		.Valid_In(bn48_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(rl48_Valid_Out)
	);
//////////KERNEL49//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110100100101100111000011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110111100111101101110101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111100000010111000000110101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111101101001101110001110000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111110101001010011101110100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111110100111000000011011111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111101101100011101001010101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111110011110011100000010000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111111011100000011100010111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111101110001001010010111011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110110010101101000100011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111101010110000110010111101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111100100111100001010010010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111111000011111000011111010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110000111011111010001001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111110100111011011110110000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111110001111010010000111011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111110101110111011000000010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110000111101100101110001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111110101001100101101110101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110001101111011101011011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111110000111111111011001001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110111011010001001111100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111110111101100010101100110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111110100111000101010111010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110000110100111010101100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111101100000010000000010110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111111100001110000101010110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111011100010001011110101000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110000001001010100100010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111110100101101010110001001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111101100101100110010001000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111110101110110100111010011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b00111110101010101000010101011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111110000011001011100000010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111111000001011010010110001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b10111110001010110010010001000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111100101010111011110111110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111101100001100010000010010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111110100101001001010100110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111110001101100110111001000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111110110001100000000010010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111111011010110011110010001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111110100010110000101010000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111110100110101111010110111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b10111110001011111101010110100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111111001010010000101111011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111110100001010100011000011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b00111101110101110000101101001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b00111101110101101111010101000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b10111111011101100010010011101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b10111100111110001011101001000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b00111110001001110001010100000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111110101101101100001000000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111110001111110100100111111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111110001011100110001101101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111110110000110111010110000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111110110111101010001101010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b10111110000101111001100111100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111111001101011111000001101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111110100101011100101101111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111111000000000010111101000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b10111110101010010101001011100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111110010010110001000001001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel49_Valid_Out)
	);
	Adder_64input add_k49(
		.Data1(Data_Out_Kernel49[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel49[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel49[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel49[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel49[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel49[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel49[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel49[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel49[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel49[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel49[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel49[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel49[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel49[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel49[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel49[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel49[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel49[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel49[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel49[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel49[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel49[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel49[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel49[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel49[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel49[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel49[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel49[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel49[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel49[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel49[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel49[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel49[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel49[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel49[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel49[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel49[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel49[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel49[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel49[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel49[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel49[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel49[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel49[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel49[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel49[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel49[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel49[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel49[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel49[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel49[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel49[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel49[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel49[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel49[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel49[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel49[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel49[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel49[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel49[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel49[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel49[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel49[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel49[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel49),
		.Data_Out(add_k49_Data_Out),
		.Valid_Out(add_kernel49_Valid_Out)
	);
	Batch_Norm bn_kernel49(
		.Data_A(32'b00111110111011100000011101011001),
		.Data_B(32'b00111111010011001011101100011010),
		.Data_In(add_k49_Data_Out),
		.Valid_In(add_kernel49_Valid_Out),
		.Data_Out(bn49_Data_Out),
		.Valid_Out(bn49_Valid_Out)
	);
	Relu_Core rl_kernel49(
		.Data_In(bn49_Data_Out),
		.Valid_In(bn49_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(rl49_Valid_Out)
	);
//////////KERNEL50//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110100001000111111000001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111111001011001000100101111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110100110010001101010110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111101011000100001100011010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111110000110000000111100100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110100100101001010011001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111110000110100110001101100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111110101001100111111000000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111100001100110101101000101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110111000111001000100011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110110001110100110110011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111101110110000100100100100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111101011111000000110101000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111110111000001111011100010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111101010111100010010010101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111010101000010010100001101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110101101100101110011101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111111000001110000101001101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111101110011111100010100101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111110100001111101010010010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111101100100001101111110000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111101111011000000011101101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111111000110011110110110011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111111011011011010110111101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111111001001001001100011110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111101101011110100100001011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111111000010010111011010100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110110100011011010101000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111111000010000111001100101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110010110001111001001111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111110110001111010000000000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111110101001111010011101110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111110101111011010011110001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111110100111111011100001110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111111000100101100111111110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111110000001000010101000000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b10111110101101110000001000001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111101000000110011111011111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b00111011111101010100100010111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b00111101010111111010011100111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b10111111001010010101100101010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b10111101110110110111011111111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111110111001011010111110011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111101101101101110100000011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b00111100011011100000000000101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b10111111000010110001010101000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b10111101010010101100110111111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111101011000100101011111100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b00111110101000111111100110001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b00111101111011111100111011000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b10111110000110010111111111111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b10111101100101000100111000101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111100001000100110111001110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111110111110100000100000101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b10111111001011011111111110101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b00111101100100110101101101110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111110011111000001100100100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111110011011000110100001100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111111000110110000011001010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b00111110010010001101011111100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111111001111011000010110111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111110111011110011101110010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111110101001011010111111111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b10111110010100111111010110000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel50_Valid_Out)
	);
	Adder_64input add_k50(
		.Data1(Data_Out_Kernel50[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel50[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel50[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel50[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel50[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel50[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel50[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel50[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel50[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel50[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel50[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel50[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel50[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel50[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel50[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel50[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel50[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel50[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel50[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel50[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel50[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel50[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel50[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel50[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel50[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel50[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel50[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel50[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel50[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel50[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel50[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel50[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel50[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel50[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel50[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel50[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel50[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel50[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel50[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel50[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel50[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel50[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel50[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel50[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel50[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel50[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel50[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel50[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel50[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel50[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel50[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel50[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel50[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel50[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel50[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel50[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel50[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel50[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel50[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel50[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel50[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel50[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel50[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel50[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel50),
		.Data_Out(add_k50_Data_Out),
		.Valid_Out(add_kernel50_Valid_Out)
	);
	Batch_Norm bn_kernel50(
		.Data_A(32'b00111110111001010010100100011110),
		.Data_B(32'b00111101000100010101100011001101),
		.Data_In(add_k50_Data_Out),
		.Valid_In(add_kernel50_Valid_Out),
		.Data_Out(bn50_Data_Out),
		.Valid_Out(bn50_Valid_Out)
	);
	Relu_Core rl_kernel50(
		.Data_In(bn50_Data_Out),
		.Valid_In(bn50_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(rl50_Valid_Out)
	);
//////////KERNEL51//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110100001000100101111010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110101110011010111101100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111111001110000000001100000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111101010010100100001000101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111110011110001011111011000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110110101110010101000110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111110101001110001101100001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111110110001101101001100101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110001111111011110100001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111011100011010110010011000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110101001011100010110110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111101110101010001011001101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111110010001100110101000011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111111010100101001000111101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110100001010110100100101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111101011101100001001111001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111100100010111011010100111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111101100000101101110000110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111011011000001100000101111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111100110110010111011101110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111111000101111110110101100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111110001110111000001010001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110010110000110100100101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111101101101001011100001000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111111000000001110100000010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111101111101000111111001101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111101110011111100100100110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110110011000000011101001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111111000011111010110100011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110110111010001011111011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111110001101001001111000100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111110001110101110001001001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111101100101110101000100110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111010010111110101110110110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111111101000100000001110000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b10111110100111011111010110010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b10111110011100010111011011111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b00111101101111011001110110111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b00111110011101111101111111111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b00111111000111110110011010000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111110100111101110111011110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111110111110111111101011100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b00111101101001001011100011001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111101110111011100100000111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111110001100000110010101111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111011001110111110111111111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b10111110110111101111110010010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111110101000011101111001010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111100000011110010011001000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b00111110101110100001001101111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111111000100011000101110100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b10111110011101000011100010100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b00111110011010110010011010101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b00111110111110100000011011100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111101001111101001100100001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111100110011111100101101101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b10111110011001000111010001010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b10111110010001000011011010010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111101110110001101100100110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b00111110111000010011110010101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b10111110100010000011101110111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111101100100010000101111011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b10111111001001011101100110010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b10111110100101011010000011110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel51_Valid_Out)
	);
	Adder_64input add_k51(
		.Data1(Data_Out_Kernel51[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel51[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel51[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel51[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel51[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel51[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel51[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel51[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel51[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel51[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel51[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel51[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel51[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel51[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel51[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel51[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel51[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel51[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel51[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel51[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel51[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel51[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel51[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel51[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel51[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel51[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel51[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel51[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel51[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel51[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel51[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel51[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel51[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel51[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel51[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel51[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel51[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel51[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel51[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel51[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel51[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel51[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel51[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel51[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel51[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel51[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel51[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel51[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel51[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel51[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel51[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel51[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel51[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel51[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel51[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel51[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel51[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel51[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel51[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel51[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel51[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel51[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel51[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel51[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel51),
		.Data_Out(add_k51_Data_Out),
		.Valid_Out(add_kernel51_Valid_Out)
	);
	Batch_Norm bn_kernel51(
		.Data_A(32'b00111110111101101110010010111101),
		.Data_B(32'b10111110011100010001010000011011),
		.Data_In(add_k51_Data_Out),
		.Valid_In(add_kernel51_Valid_Out),
		.Data_Out(bn51_Data_Out),
		.Valid_Out(bn51_Valid_Out)
	);
	Relu_Core rl_kernel51(
		.Data_In(bn51_Data_Out),
		.Valid_In(bn51_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(rl51_Valid_Out)
	);
//////////KERNEL52//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111101011000001000101001011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111111000010010111101001100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111111000010101101001001100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110011101010101001100001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111111000011001111000001001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111101100100100000100011111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111101101101101100001000011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111110110110110110001000001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110111101101100101001111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110110111011100010100000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110101011011010111111001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110111010111000111001011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110111110011010101010010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111101010111000011110100101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111101101110011111100100000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111110011110100000001000111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110000010110110100101010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111111000001010101001110000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111101110000100000000001000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110000110111110010010110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110011011101101100101111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111110000011101111101011010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111101100100101100101100110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111110011000101100111001100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111110100100010111001100001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110010110110110000011010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111111000100110000100001001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111101100110011011100111111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111110100010111010100000100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111111001110100000011000101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111101111001111110001111110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111111010000000000111010101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b00111110101111001011110111001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111111010010101110111010110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111111000000010010001100100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111101001110000101010001010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111110000110011111001011110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b00111110001000110010111000100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b00111110101100100110011111000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b00111110101001010000000101110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b10111100111100101100000110001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111110111001000101000110111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b00111111000001011101010100010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b00111110010010101000011001111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111110101110111100110000101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b10111110001110001011110000110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b10111110001000010011100010100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111111000000100110000111111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b00111111001101001000111110101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111110111000001111001000100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b10111110010101010001011000000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b10111110100111011000011010010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b00111110100110101111001110001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b00111101101101111111010100011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b10111101110010001110101000101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111111010010110101000010000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111110010010101000100000101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111110001110110011101001000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111101110000011111010110110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b00111100110000010011000110011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b10111110111001000111101010111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b10111100110111111110111110100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b10111101011100100000100011000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111110100110010100010100100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel52_Valid_Out)
	);
	Adder_64input add_k52(
		.Data1(Data_Out_Kernel52[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel52[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel52[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel52[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel52[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel52[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel52[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel52[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel52[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel52[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel52[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel52[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel52[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel52[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel52[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel52[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel52[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel52[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel52[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel52[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel52[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel52[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel52[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel52[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel52[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel52[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel52[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel52[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel52[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel52[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel52[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel52[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel52[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel52[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel52[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel52[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel52[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel52[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel52[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel52[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel52[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel52[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel52[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel52[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel52[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel52[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel52[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel52[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel52[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel52[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel52[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel52[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel52[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel52[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel52[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel52[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel52[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel52[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel52[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel52[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel52[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel52[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel52[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel52[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel52),
		.Data_Out(add_k52_Data_Out),
		.Valid_Out(add_kernel52_Valid_Out)
	);
	Batch_Norm bn_kernel52(
		.Data_A(32'b00111110101111000001110000100001),
		.Data_B(32'b00111111001110001011111110000011),
		.Data_In(add_k52_Data_Out),
		.Valid_In(add_kernel52_Valid_Out),
		.Data_Out(bn52_Data_Out),
		.Valid_Out(bn52_Valid_Out)
	);
	Relu_Core rl_kernel52(
		.Data_In(bn52_Data_Out),
		.Valid_In(bn52_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(rl52_Valid_Out)
	);
//////////KERNEL53//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110111000100001111100001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111110011101100010111100100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110001100011111111110010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110101101011101101001011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111111001001110000000110101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111110101011011011111010100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111101101010111101100100111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111110111010011101110110011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110001000011111010101101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110100110101100001110011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111110100001101110110000110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111110000101100010010010110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110100011011110011110000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111110001100001101001000100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111111000010110001001010100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111110001100111110010000100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110100011101001010000100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110010101010101111001100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111111001101100001001010011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111101101011111111111111011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110100000010001110011010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111100011110100100000110001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111111000011000111100101001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111101010110000011010010011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111110101101010111101101111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110011110100001010001001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111110101001100010011101001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110100011101001111100110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111111001101001000000010110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111110110110110101000011000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111111001000000110010111111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111111001001011111100001110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111111000110000010110101111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b00111111000101001000011110110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111110101011111110111110100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111011100101010011001100111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b10111110110001011100000100000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111011101101011001111110000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111110000001101001110010000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b00111110011000010000001110010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b10111111010000011000011011101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b10111110110011011100011000101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111101100110100101001010011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b00111110001100010111110010010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111101110001110110111101010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111110110100101101001101000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b10111110100001000011101110110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b00111110111011000110110100011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b00111111000100010101001100011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b00111101000100111110100001011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111110110100100111001101010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111111000110001100101101100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111101100101101000001010010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111110011010101111101100011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b10111110100101111011000111101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111110110101010110101011100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111110110000101011110110010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111101101001011110101100110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111110010101101010001100000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b00111110001110010000101110001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b10111110101010101011000100010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111110100111111110100100000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111110100011101111011001101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111011110110011001011110001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel53_Valid_Out)
	);
	Adder_64input add_k53(
		.Data1(Data_Out_Kernel53[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel53[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel53[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel53[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel53[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel53[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel53[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel53[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel53[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel53[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel53[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel53[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel53[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel53[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel53[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel53[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel53[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel53[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel53[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel53[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel53[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel53[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel53[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel53[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel53[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel53[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel53[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel53[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel53[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel53[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel53[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel53[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel53[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel53[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel53[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel53[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel53[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel53[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel53[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel53[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel53[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel53[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel53[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel53[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel53[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel53[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel53[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel53[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel53[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel53[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel53[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel53[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel53[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel53[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel53[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel53[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel53[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel53[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel53[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel53[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel53[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel53[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel53[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel53[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel53),
		.Data_Out(add_k53_Data_Out),
		.Valid_Out(add_kernel53_Valid_Out)
	);
	Batch_Norm bn_kernel53(
		.Data_A(32'b00111110111100110011111001110000),
		.Data_B(32'b00111111000011101110110001000000),
		.Data_In(add_k53_Data_Out),
		.Valid_In(add_kernel53_Valid_Out),
		.Data_Out(bn53_Data_Out),
		.Valid_Out(bn53_Valid_Out)
	);
	Relu_Core rl_kernel53(
		.Data_In(bn53_Data_Out),
		.Valid_In(bn53_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(rl53_Valid_Out)
	);
//////////KERNEL54//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110101110000010001110001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111110000100010011000110011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110100100101011110001001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110110011000001001000111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111110111110101101000100100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111111001000111110011100001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111100110011100101001100000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111110100101001101110010010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111101010010110000011110100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111111001111001101011111111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111110110011000111111001011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110101001100001000110011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111101111000101010001010100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111110101011010001101110100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110001011011100110100110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111110010011000111100110110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111101100101011111110100001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110101000010010111100001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111101100110101101011011001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111101010000010111110010100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110000111010111000101001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111110110100111101111010100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110110100100110101100011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111110110011000011110010101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111110010000110001111111110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111111000100110000101101000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111101101110100000011010110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111110100111101101010101010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111110111101000111010001000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111110010111101110010011110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111101111001100010110000001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110010010101100011010011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b00111110101001001100110001000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111110110011001111101100001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111100011111110110110101001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111110001000100001111000011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b10111110000110000010001101010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111100101110111111010110011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111110111001011011110000001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111111000011000110101110011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b10111101110011001001100000010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111110011111000100000001011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111110110110001110101000111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b00111110110100111010010000011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111110000011010111011001011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b10111110000111111111001001110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111101000110000001000100101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b00111110110101110000111010000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111100100111010110011000010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b00111100001100011001101111010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111111000100010110010110001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111110110010110000011011001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111110111101111101000100001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111110100000000101110110010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b10111111010101011101100110101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b00111110010010110111101111110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111110001111011110010010001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111110110101101010111001001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b10111101111100011100000000010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b00111111000110011101101010000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111111000000100001100101011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111100111110001001111100110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b10111110101010000000110011100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b10111110011010001001010000011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel54_Valid_Out)
	);
	Adder_64input add_k54(
		.Data1(Data_Out_Kernel54[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel54[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel54[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel54[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel54[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel54[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel54[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel54[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel54[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel54[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel54[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel54[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel54[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel54[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel54[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel54[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel54[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel54[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel54[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel54[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel54[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel54[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel54[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel54[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel54[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel54[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel54[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel54[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel54[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel54[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel54[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel54[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel54[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel54[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel54[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel54[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel54[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel54[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel54[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel54[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel54[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel54[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel54[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel54[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel54[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel54[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel54[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel54[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel54[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel54[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel54[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel54[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel54[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel54[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel54[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel54[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel54[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel54[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel54[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel54[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel54[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel54[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel54[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel54[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel54),
		.Data_Out(add_k54_Data_Out),
		.Valid_Out(add_kernel54_Valid_Out)
	);
	Batch_Norm bn_kernel54(
		.Data_A(32'b00111110111100001000100011001011),
		.Data_B(32'b10111111000111101001110100101111),
		.Data_In(add_k54_Data_Out),
		.Valid_In(add_kernel54_Valid_Out),
		.Data_Out(bn54_Data_Out),
		.Valid_Out(bn54_Valid_Out)
	);
	Relu_Core rl_kernel54(
		.Data_In(bn54_Data_Out),
		.Valid_In(bn54_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(rl54_Valid_Out)
	);
//////////KERNEL55//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111111000011100100100000000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111110101000010000000110010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111111000000000001100001110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110100101111100101101101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111110000100111010001010111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111101100110100011101011101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111110110100011010100110001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111110010011000101101111101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111110101111101101000000110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111110100101001011101001011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110110000110011100001101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110000111011000011011000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111101010111001100011011011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111101110011100010001000000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111111010101011101010110001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111111000000101110110111101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111110101100010001110111011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111101110111000001101010001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110100110111010011010100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111101000101000111100111010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111111000100000101111000111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111111000000111111011110111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111101100010111101011111111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111111000101010101010100110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111111000100111111000000010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110111100000111010100000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111111000000101010101111011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110000011001111000010111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111110111001101011010011100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110000110110001001000010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111100011010111100001011111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110101100000100001001110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b00111110100100111010001101111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111110001100011011100010101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111111001011100001011000011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b10111110100010001000001101000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b10111110100100011100100110001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111110111011010011000010000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111110101111111010011010001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b00111110010000011101000111110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b10111110100011011011110101000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b10111110100000101001100100010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b00111110100011100111100100101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111111000110000001011010110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b00111110010001100011101110000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111101010000110011001010100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b10111110111010110010111100100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b00111110110010111001100011110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b00111100010110011001100110101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b00111101111100000100100000101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b10111110100001100010001000100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111110100100011101001000100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111110000111100010111001010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b00111100111011100010111010111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b10111110101110110101001111000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111111001001101111111101111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b10111110011010010010000110100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111101110111000111100011110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b10111110000011000011111010000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b00111110101001110101111101001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111110110000111111011100100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111110110110001100001010001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111110100110111110010011001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111111001011010011010111100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel55_Valid_Out)
	);
	Adder_64input add_k55(
		.Data1(Data_Out_Kernel55[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel55[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel55[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel55[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel55[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel55[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel55[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel55[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel55[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel55[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel55[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel55[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel55[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel55[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel55[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel55[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel55[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel55[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel55[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel55[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel55[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel55[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel55[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel55[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel55[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel55[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel55[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel55[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel55[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel55[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel55[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel55[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel55[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel55[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel55[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel55[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel55[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel55[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel55[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel55[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel55[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel55[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel55[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel55[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel55[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel55[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel55[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel55[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel55[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel55[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel55[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel55[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel55[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel55[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel55[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel55[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel55[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel55[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel55[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel55[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel55[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel55[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel55[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel55[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel55),
		.Data_Out(add_k55_Data_Out),
		.Valid_Out(add_kernel55_Valid_Out)
	);
	Batch_Norm bn_kernel55(
		.Data_A(32'b00111110110111111111110100010100),
		.Data_B(32'b10111101001111001000010010100000),
		.Data_In(add_k55_Data_Out),
		.Valid_In(add_kernel55_Valid_Out),
		.Data_Out(bn55_Data_Out),
		.Valid_Out(bn55_Valid_Out)
	);
	Relu_Core rl_kernel55(
		.Data_In(bn55_Data_Out),
		.Valid_In(bn55_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(rl55_Valid_Out)
	);
//////////KERNEL56//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111110100110101101100100101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111110110001011111101111011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110111010001110001011100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110101010100101010110101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111101100110000011000010010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111110100001101110011100100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111000101110001010010010100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111101100001111100111010111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110000110000110101101111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110010011001001100110011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110000101110011111101110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111111001100001011101011101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111110000011001011001100100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111110111001011001111010110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110011001100000101011010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111111011111010111111011010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110011100001100011010010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111100100111100010000011101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110011010000000010000110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111101101111110010011100000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111101101100011111100011101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111101100000000011000110101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110001000111111000100001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111110001111111011001010010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111110010010001110000100111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111110010011000110101010011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110100000001111010011101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110100010100100111111101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111110000001111111100110110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111101110100001110000100111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111110001000111110100011010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110101000000001010010111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111110011101110110011110111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111111001000111100100101101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111111000010101100101110011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111110100100001101101111000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b10111101100000100100010100011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b00111110000110101111101111000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b00111110101011010010110101010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b00111101101010011101010100101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111101100101111111100101001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111111000011001100100000101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111110001100100011111011000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111100111010011010000001010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111110100010000000111011101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b10111111010101000011100100111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111110101101101000011010111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b00111110110110110000001001101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b00111111001100101100001100011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111110001111100001111000000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111111000001010100001010011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b10111110111000011010010000101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111110110101110001110111000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b00111101100100011001001101001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111111000100010111001110110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111110110000111011111110000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111100111110011010011001110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111101110011010011101101011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b10111110101011110001101101100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111110101101010011001001110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b10111110011110110000101001011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111110110011110001101111010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111101010110100101100100100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111110010101011001001010111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel56_Valid_Out)
	);
	Adder_64input add_k56(
		.Data1(Data_Out_Kernel56[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel56[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel56[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel56[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel56[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel56[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel56[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel56[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel56[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel56[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel56[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel56[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel56[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel56[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel56[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel56[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel56[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel56[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel56[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel56[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel56[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel56[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel56[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel56[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel56[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel56[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel56[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel56[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel56[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel56[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel56[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel56[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel56[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel56[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel56[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel56[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel56[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel56[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel56[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel56[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel56[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel56[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel56[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel56[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel56[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel56[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel56[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel56[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel56[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel56[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel56[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel56[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel56[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel56[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel56[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel56[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel56[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel56[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel56[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel56[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel56[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel56[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel56[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel56[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel56),
		.Data_Out(add_k56_Data_Out),
		.Valid_Out(add_kernel56_Valid_Out)
	);
	Batch_Norm bn_kernel56(
		.Data_A(32'b00111110111011011001000000010100),
		.Data_B(32'b00111100101011010011101100101111),
		.Data_In(add_k56_Data_Out),
		.Valid_In(add_kernel56_Valid_Out),
		.Data_Out(bn56_Data_Out),
		.Valid_Out(bn56_Valid_Out)
	);
	Relu_Core rl_kernel56(
		.Data_In(bn56_Data_Out),
		.Valid_In(bn56_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(rl56_Valid_Out)
	);
//////////KERNEL57//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110001111100000100110000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111110001101110000000101111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110101101010000000100011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111111000111111111011000011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111110110111100101101110001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110110100011000101000110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111110100001010100111011000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111110100100100100101101101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111100100011100000101111010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110111110111100010001000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111011101110000011001111001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110000001110001011000000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111111000000011011011001111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111110100001100100100101101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110000011100100001001010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111111001010010010101110101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111110100100100100101111100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111110100111111000010001000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110011101101101110101110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111111101001010000000101000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111101001100001000001101101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111100000010011110001000010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110101010110111001001010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111110111101011000000100110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111011011111001100101100101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111100101111001111110100010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111111000101101001111100100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111100100000100101001100011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111110101101001000101000001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110101000110010010100100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111110000101011001000011101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111101110110110000000110011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b00111101110110001100000011011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111111011010011000101011010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111110011100101001111001110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111110001101101100101100001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b10111110101110100110010001011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111110011110110011100101110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b00111110000011111011010010110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b00111110101001111111000110110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111110101011101110100111000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b10111110100001011110000000010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b00111110010011100101101000010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b00111110101000111110000111110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111111000010001110011010110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b10111100101100111001000011110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111110110000111100101010111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111110011010001011101110101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b00111111100000111001010101110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b00111101011001000100011111010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111110001100101001011100101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b10111110111001100100011111000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b00111110000110101010001100111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b00111101100101110110111010111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111110000001011010100011101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111110001001100010101000101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111110000011000001000100100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111110010001010000101010110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111100010011100001000110011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b00111110011001000110100100000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111110111010000001111111001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111111000000000100010011011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b10111100111000001110001100111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b10111101000101101011100100010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel57_Valid_Out)
	);
	Adder_64input add_k57(
		.Data1(Data_Out_Kernel57[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel57[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel57[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel57[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel57[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel57[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel57[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel57[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel57[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel57[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel57[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel57[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel57[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel57[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel57[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel57[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel57[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel57[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel57[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel57[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel57[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel57[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel57[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel57[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel57[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel57[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel57[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel57[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel57[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel57[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel57[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel57[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel57[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel57[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel57[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel57[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel57[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel57[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel57[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel57[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel57[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel57[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel57[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel57[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel57[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel57[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel57[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel57[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel57[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel57[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel57[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel57[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel57[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel57[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel57[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel57[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel57[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel57[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel57[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel57[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel57[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel57[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel57[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel57[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel57),
		.Data_Out(add_k57_Data_Out),
		.Valid_Out(add_kernel57_Valid_Out)
	);
	Batch_Norm bn_kernel57(
		.Data_A(32'b00111110110010001001011111001001),
		.Data_B(32'b00111110111101100000010101101011),
		.Data_In(add_k57_Data_Out),
		.Valid_In(add_kernel57_Valid_Out),
		.Data_Out(bn57_Data_Out),
		.Valid_Out(bn57_Valid_Out)
	);
	Relu_Core rl_kernel57(
		.Data_In(bn57_Data_Out),
		.Valid_In(bn57_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(rl57_Valid_Out)
	);
//////////KERNEL58//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110100100000011110101010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110100101110001110000010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111111000100001010011100011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110101001100010001011111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111110110010010011110001100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111111000011111101100110001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111110001110101110100000000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111110101001110101100100100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111110010010100010101001100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111111001100011101001111001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111110111111000110101100100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111101001100110010010100101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111110111010010000101100001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111110011100101101100101000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110101010101001111001111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111100000101100100110110100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110100100011111110111000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111110010111000111010101001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111100000110111100110100111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111101000111110101011100010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111111100110001011100011100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111101100011110010000111000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111101101000101111000110011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111111001100110000111110011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111110100111110000110110111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110010010011011100101010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110001101000010111100010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111110100100000010110000000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111110001001001101000111110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111111000010101001011110010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111110011101100110000110011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110001110000011010111101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b00111110110000101100000100100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111110101110001110011010001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111110101000110000100001111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111110101001101100010001101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111101000001111000001101000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b00111110110111110100010110100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b00111110101001011110101100010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111111000001011011111100000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b10111100111010011100111000011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111100101100010111110011110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111101111011011001000100010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b00111110111101011000110010101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b00111101101101101000001000111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b10111110100010001000011101001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b10111101110111011010000110100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111111000000010010111010110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b00111110100011110010101110111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111110101111010011011101111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b10111110101000000010001001110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111101111011111010001100111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b00111111011001011001101100000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b00111101000100001010111100100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b10111110001011110011101001111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111110110001001001100011100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b10111110110100110011110001010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b10111111000000100000001000110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111110010011000111001110111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111110110101011000111100110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b10111100101111110111010101001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b10111110111001100010000001110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111110100101110010010110111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111110111101010010100100000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel58_Valid_Out)
	);
	Adder_64input add_k58(
		.Data1(Data_Out_Kernel58[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel58[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel58[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel58[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel58[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel58[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel58[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel58[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel58[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel58[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel58[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel58[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel58[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel58[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel58[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel58[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel58[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel58[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel58[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel58[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel58[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel58[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel58[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel58[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel58[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel58[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel58[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel58[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel58[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel58[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel58[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel58[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel58[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel58[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel58[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel58[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel58[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel58[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel58[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel58[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel58[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel58[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel58[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel58[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel58[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel58[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel58[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel58[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel58[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel58[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel58[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel58[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel58[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel58[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel58[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel58[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel58[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel58[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel58[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel58[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel58[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel58[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel58[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel58[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel58),
		.Data_Out(add_k58_Data_Out),
		.Valid_Out(add_kernel58_Valid_Out)
	);
	Batch_Norm bn_kernel58(
		.Data_A(32'b00111110111000110001001101001110),
		.Data_B(32'b00111111000000101000101111111001),
		.Data_In(add_k58_Data_Out),
		.Valid_In(add_kernel58_Valid_Out),
		.Data_Out(bn58_Data_Out),
		.Valid_Out(bn58_Valid_Out)
	);
	Relu_Core rl_kernel58(
		.Data_In(bn58_Data_Out),
		.Valid_In(bn58_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(rl58_Valid_Out)
	);
//////////KERNEL59//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111011010011101101011100100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111101101010011011001000010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110100111000110001000010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110001111000111001000111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111111000001111110101010101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110100000111000110111011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111111000001101011000001011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111110101010011011101100100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110100111010010101111001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111101101010110001000110010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111110100000101010101111000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111111000001110010000110100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110100110001111001011011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111110101100010011110011010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111111011011111111100100000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111110001010010110100010010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111110101001000000101000000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110101010011001001011000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111101110001000010101110010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111011001100011110101010101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111101111000100000100001111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111110100111101100010101111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111110000010010111010011101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111110011000011000000001001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111111000100111011100111001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111101110101000111010000011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110101010010111100111111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111110011100101011001100101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111110110100011011011000010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111111001111011110011000101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111101000010000001010001010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110011011100110001010011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b00111101100110101110101110001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b00111101001110100010010111000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111110101110001010100101110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b10111110111001110101101000100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b10111110000001001011010111001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111110110000000100110101110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111110111111101001010111000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b00111110111101011100011100100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b10111110011001111001011110101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b10111101111001000111001101110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b00111110101100101101111101011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b00111110011111011101001010100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111110100101010111101000010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111111011010000111011111000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b10111110110110100110100110010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111110001100111011110110110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b00111110101011011000111010101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111101011000110110000101100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b10111011011011000101101111100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111111000001010000100100110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111110010011011001100000000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b00111101011100010000110001001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b10111111010001011000001111010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111101011000011011001001101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111110000101001010000110001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111110110010000010001101100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111101101010101001101101101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111110010001111110111010000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111111000011111100111011000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111110101101010100101101011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b10111110000010000110101010001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b10111111000111000111110111110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel59_Valid_Out)
	);
	Adder_64input add_k59(
		.Data1(Data_Out_Kernel59[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel59[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel59[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel59[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel59[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel59[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel59[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel59[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel59[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel59[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel59[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel59[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel59[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel59[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel59[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel59[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel59[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel59[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel59[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel59[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel59[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel59[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel59[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel59[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel59[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel59[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel59[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel59[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel59[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel59[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel59[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel59[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel59[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel59[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel59[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel59[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel59[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel59[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel59[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel59[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel59[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel59[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel59[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel59[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel59[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel59[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel59[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel59[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel59[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel59[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel59[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel59[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel59[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel59[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel59[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel59[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel59[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel59[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel59[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel59[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel59[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel59[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel59[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel59[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel59),
		.Data_Out(add_k59_Data_Out),
		.Valid_Out(add_kernel59_Valid_Out)
	);
	Batch_Norm bn_kernel59(
		.Data_A(32'b00111110111000001011111100010101),
		.Data_B(32'b10111101110001110011011100000001),
		.Data_In(add_k59_Data_Out),
		.Valid_In(add_kernel59_Valid_Out),
		.Data_Out(bn59_Data_Out),
		.Valid_Out(bn59_Valid_Out)
	);
	Relu_Core rl_kernel59(
		.Data_In(bn59_Data_Out),
		.Valid_In(bn59_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(rl59_Valid_Out)
	);
//////////KERNEL60//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111100111101110101011101101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111100010001101111111000110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110000000010110011010101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110000101000010110010001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111101101010010000001000111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111101101100100000110100110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111110110100010000001100100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111111001010010010000010000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111100110010000001110100100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111110100111110010011001000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111101110010011110100110100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110010100000111010000000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110101100100000011110000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111101110001101110110011111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110111011101010100011100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111110001010000011001000000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110000101001010101110010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111111101011010110111001101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110110101100101000011111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111101111010111010100111100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111101110100110111110000101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111111000101101000110011011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111100000001011101111010100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111111000001001011000010111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111101001101101111001001001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111111001100001001110010111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111101101000110000100111101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111110011001001000011010001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111110011010111010010100100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111111011010011001101000010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111110000101110000001101011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110000111000000011001010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111111000000100001100001011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111110100001111010110000100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111111000101000110010000100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b10111110101001110011100010011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b10111101101010111100001101000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111101111110101010011010001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b00111110000010101011000010100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b00111110101011100000101100100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111100100100101001001111101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b10111111001011000110110000001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111101101000101110101000100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111110001011101110001010101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b00111101111110011010110110111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111110011010110001011110011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b10111101101111100111101111001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111110110001110000001100100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b00111110101001001110101001110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111110110111101000001110010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b10111101001111001001101100110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111110111010110101110101101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b00111110111010011010010111110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b00111101101100111001010011111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111110101001011111111111000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b00111011110110110110100101101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b10111110111110110010100011110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111110110010100010110011100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111110000001001100110001100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b00111111000011010011010111000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111110001001010110010010110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111110010101101011110010110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b10111110101101000001010110110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b10111110100100011110100000110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel60_Valid_Out)
	);
	Adder_64input add_k60(
		.Data1(Data_Out_Kernel60[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel60[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel60[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel60[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel60[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel60[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel60[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel60[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel60[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel60[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel60[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel60[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel60[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel60[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel60[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel60[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel60[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel60[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel60[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel60[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel60[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel60[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel60[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel60[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel60[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel60[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel60[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel60[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel60[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel60[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel60[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel60[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel60[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel60[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel60[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel60[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel60[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel60[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel60[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel60[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel60[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel60[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel60[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel60[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel60[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel60[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel60[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel60[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel60[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel60[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel60[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel60[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel60[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel60[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel60[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel60[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel60[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel60[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel60[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel60[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel60[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel60[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel60[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel60[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel60),
		.Data_Out(add_k60_Data_Out),
		.Valid_Out(add_kernel60_Valid_Out)
	);
	Batch_Norm bn_kernel60(
		.Data_A(32'b00111110111100011110011000101010),
		.Data_B(32'b00111111001100100011101100111100),
		.Data_In(add_k60_Data_Out),
		.Valid_In(add_kernel60_Valid_Out),
		.Data_Out(bn60_Data_Out),
		.Valid_Out(bn60_Valid_Out)
	);
	Relu_Core rl_kernel60(
		.Data_In(bn60_Data_Out),
		.Valid_In(bn60_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(rl60_Valid_Out)
	);
//////////KERNEL61//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111110100000100011011111010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111111000010011010010101010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111010110001010010100100010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110110101100101000100100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111110111101011100101110101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111110010010111111000001000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111110101000010111000001100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111101000011001111100000111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110100111000000000111101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111101101001011100010001000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111111000000001011001111000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111101110001001111000101011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111111010101010110000110000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111101000011100010100000010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111101101111011010111111111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111111010111010000000110001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111110110100110101010101000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111111000100100101011000111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111110011001100110101001000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111110001110110101110110100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110001010101001011100110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111110100010110110000110001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111111000101010111100100101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111101110110011000110011100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111110110110001010000010100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111101111010101001000101110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111110011110101011100101011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111111001111101010000110010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111101010010101110110110111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111110100101000010100011000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111110111001011011100101100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110011010011000000000101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b00111111001110011101101101000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111111001101110011000110110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111110101000100101111110011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111111000010001111110110010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b10111110100101100011110101110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111110010000001100101111100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111110101000111111001001001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111110001010011110000001110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111110111000001101110111001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b10111100111001110010101011111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b00111110100100111010010100101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111110101000110110011110010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111101100000011010000100010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111101110001110101100110110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b10111101110000101000001001011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b00111110001110110011011011010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111110000001101110000100110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111110101100000110101111010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111110101010111011100010111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111110110101101101000101111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b00111110010111101100011111110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b00111110000110010100100111001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b10111101100101000011110111101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111111000100101000010110011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111101111110001011100110111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b10111101110001100100100011110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b10111110111011011100001110111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b00111110101111000110100111000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b10111110100011101110001111101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b10111110010000001100100000001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111111000101011011000100010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111110100011111011001000100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel61_Valid_Out)
	);
	Adder_64input add_k61(
		.Data1(Data_Out_Kernel61[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel61[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel61[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel61[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel61[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel61[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel61[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel61[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel61[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel61[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel61[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel61[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel61[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel61[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel61[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel61[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel61[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel61[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel61[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel61[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel61[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel61[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel61[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel61[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel61[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel61[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel61[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel61[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel61[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel61[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel61[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel61[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel61[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel61[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel61[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel61[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel61[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel61[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel61[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel61[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel61[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel61[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel61[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel61[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel61[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel61[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel61[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel61[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel61[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel61[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel61[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel61[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel61[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel61[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel61[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel61[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel61[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel61[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel61[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel61[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel61[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel61[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel61[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel61[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel61),
		.Data_Out(add_k61_Data_Out),
		.Valid_Out(add_kernel61_Valid_Out)
	);
	Batch_Norm bn_kernel61(
		.Data_A(32'b00111110110100110100001110001111),
		.Data_B(32'b00111111100111111011000100111001),
		.Data_In(add_k61_Data_Out),
		.Valid_In(add_kernel61_Valid_Out),
		.Data_Out(bn61_Data_Out),
		.Valid_Out(bn61_Valid_Out)
	);
	Relu_Core rl_kernel61(
		.Data_In(bn61_Data_Out),
		.Valid_In(bn61_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(rl61_Valid_Out)
	);
//////////KERNEL62//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111111000010101010001110011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111111000011101100101101000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111111001111100000010110110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110011000100000001111000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111101110100100110110010011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111100100001110101000011001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111101011010000100101100101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111011101101011001000011001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111111001010010110000011011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111110000001100100010010001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110011101100111010100010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110111100111010111101011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110110011110100000001100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111100011010111010101011101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111101100010001111100101011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111110100001000001100001110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111011100100110101010100011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111110110100010011000010011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111110101000001110001110011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110001111101111010100110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111111011110011110011100000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111101000101001011010101000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111110000010100110101000001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111110111111000111010001001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111111000101011100110000100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111110110101011000100001000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111111000110100100011100100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110110101100000011101110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111110001100001000100111111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111110111101001111010101110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111110101111100010100010001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110000010001011010100110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b00111111001001001100010000000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111110010011000000101111111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111110010111000010011011110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b10111101001000111100010111000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b10111101100000000110000010101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b00111110010101011111101101111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b00111110000010111111100001000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b00111111000001010111000101000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b10111110110001000000010011110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b10111110100111101001100111110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111101000000110000100010000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111110101001101101011100111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111110100000001111101001111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111101011100110111110011001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b10111111001011011010110110011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111100000101100000110011000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b00111110110010010011101110111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111110101110110001100011011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111111000011110110010011111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111110111100001100111011010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b00111110001101101011000001100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b00111110000100001010000001101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b10111110111000010001000000001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b00111110010010010000100001010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b10111110010000101001000101001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b10111110011000110110000100000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b10111110100111011001101000111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b00111110011010110111101001010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b10111111000100000010110111101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b10111101010101101110010100011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111100110110000101010110111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111110000001000011100011001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel62_Valid_Out)
	);
	Adder_64input add_k62(
		.Data1(Data_Out_Kernel62[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel62[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel62[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel62[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel62[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel62[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel62[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel62[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel62[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel62[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel62[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel62[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel62[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel62[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel62[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel62[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel62[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel62[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel62[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel62[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel62[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel62[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel62[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel62[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel62[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel62[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel62[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel62[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel62[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel62[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel62[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel62[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel62[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel62[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel62[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel62[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel62[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel62[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel62[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel62[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel62[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel62[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel62[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel62[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel62[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel62[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel62[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel62[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel62[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel62[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel62[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel62[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel62[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel62[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel62[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel62[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel62[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel62[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel62[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel62[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel62[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel62[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel62[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel62[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel62),
		.Data_Out(add_k62_Data_Out),
		.Valid_Out(add_kernel62_Valid_Out)
	);
	Batch_Norm bn_kernel62(
		.Data_A(32'b00111110110101001110001000000101),
		.Data_B(32'b00111110100000101011101111110100),
		.Data_In(add_k62_Data_Out),
		.Valid_In(add_kernel62_Valid_Out),
		.Data_Out(bn62_Data_Out),
		.Valid_Out(bn62_Valid_Out)
	);
	Relu_Core rl_kernel62(
		.Data_In(bn62_Data_Out),
		.Valid_In(bn62_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(rl62_Valid_Out)
	);
//////////KERNEL63//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110010110000010001010011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111110000111100010110010001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110011110010001111111011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111100110111111010100000011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111110110110010101101000101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110011001011000000000000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111101010000111100100110010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111110110000010111110110101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110101111011101101101111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111110010000100111100000001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110101000101010101100110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111110100000111010111011110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111110001010110010101011000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111110000100010010101101100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111111000111111100010000100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111110101101100110111000011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111110111110011001101000001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111010100101111100110100001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111111011011010110010101111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111111000001110101111100111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111100101011010010110100100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111110101111100011111000000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110000001100111111010111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111111001101000010011110100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111110000110111011101010011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111101111001001011111110111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110100101011001001000011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111101101011000110001001011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111110000110011010001110111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111110001101000011011000001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111110110100101111101010111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110001101100111010110001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111110100101100101000110100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111110011011110100001101110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111011110100100110011010100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b10111110101101110101010010111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111111010001111110100011011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b00111101100101111010101001110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111110101011101001100110111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111111011110011110101100101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111101110000011011101000110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111111000111100011010001010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b00111101001010100000111111101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b00111101001101010111100001110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b00111100101001101101000000011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111110101111100101100111011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b10111111001111110011100100101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b00111110111001100100111001101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111100101100101111110111110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b00111101110001100010110010111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b10111110111100001100011001011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b10111110101001001111111011010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b00111110010000101100010111111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111101110110001101001010110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111101100001011010111001011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111111001011011111100010000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b10111101101101101011010001101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b10111110101101111011001101001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111100110011101111010010100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111100111101111100011010100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111110100010010100010001100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b10111110001011000111010110011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111110100010011110001010000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111110100110110011000001110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel63_Valid_Out)
	);
	Adder_64input add_k63(
		.Data1(Data_Out_Kernel63[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel63[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel63[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel63[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel63[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel63[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel63[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel63[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel63[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel63[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel63[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel63[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel63[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel63[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel63[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel63[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel63[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel63[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel63[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel63[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel63[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel63[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel63[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel63[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel63[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel63[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel63[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel63[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel63[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel63[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel63[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel63[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel63[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel63[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel63[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel63[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel63[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel63[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel63[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel63[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel63[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel63[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel63[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel63[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel63[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel63[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel63[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel63[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel63[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel63[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel63[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel63[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel63[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel63[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel63[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel63[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel63[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel63[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel63[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel63[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel63[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel63[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel63[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel63[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel63),
		.Data_Out(add_k63_Data_Out),
		.Valid_Out(add_kernel63_Valid_Out)
	);
	Batch_Norm bn_kernel63(
		.Data_A(32'b00111110110110101110111011101111),
		.Data_B(32'b00111110010001110011110111100010),
		.Data_In(add_k63_Data_Out),
		.Valid_In(add_kernel63_Valid_Out),
		.Data_Out(bn63_Data_Out),
		.Valid_Out(bn63_Valid_Out)
	);
	Relu_Core rl_kernel63(
		.Data_In(bn63_Data_Out),
		.Valid_In(bn63_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(rl63_Valid_Out)
	);
//////////KERNEL64//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111101100001001011001110101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110001001100111101001111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110101011110111100010010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110100010010100011001001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111111001101011000110111110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110011111110000000101000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111110001000110000010111101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111110100001110111001011000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110100111101101000110110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111111010100011110100001001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110011101111100010011111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111111001111111100110101110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111111011001101010100110001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111110010111111101100100111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110100100110110111111110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111110101000011010100000110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111100111101010101010110111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110110101010100111101111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111100000000110000110101010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111110100010110001011101110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111101000010001010010101001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111110110111110001101001110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111111001001001001010100100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111110100010100110111000001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111101010001001110110111010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111011010010101000111101001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110010010000101001001011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111100101001010111011111101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111101101011110001100000000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110010011001001111100101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111101000111100111111011000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111110101110110000010011011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b00111110001001010101010000100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b00111101010110011110100011011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111110101110001111000001100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111110011100010010001100111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b10111110110110100011011010111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111110101111110100110110100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111111011001111000011001110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111101100101100111010111011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b10111110100000001011111110000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b10111110110011001110011111111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111110010110010010000000011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b00111101101100010011101100001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111111001111110110010111111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b10111110110000100100001101100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b10111101100001110100011111111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b00111110100000100011000111001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b00111110001001010111010110110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111101000101110010011100101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b10111110011111101011100101111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b10111110101100000101010100100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b00111111001101001011000111100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111110100000100100101101101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b10111111001001100000011010100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111110001011000010010000100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b10111110010111010101001111011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111111000000100101101010001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b10111101000000111111111011101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111111000001001110110011110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b10111110010111011011011010100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b10111110101111011011111100101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111100101001010010101010010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111110001000001111110011110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel64_Valid_Out)
	);
	Adder_64input add_k64(
		.Data1(Data_Out_Kernel64[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel64[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel64[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel64[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel64[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel64[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel64[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel64[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel64[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel64[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel64[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel64[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel64[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel64[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel64[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel64[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel64[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel64[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel64[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel64[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel64[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel64[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel64[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel64[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel64[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel64[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel64[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel64[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel64[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel64[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel64[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel64[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel64[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel64[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel64[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel64[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel64[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel64[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel64[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel64[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel64[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel64[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel64[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel64[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel64[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel64[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel64[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel64[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel64[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel64[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel64[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel64[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel64[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel64[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel64[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel64[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel64[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel64[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel64[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel64[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel64[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel64[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel64[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel64[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel64),
		.Data_Out(add_k64_Data_Out),
		.Valid_Out(add_kernel64_Valid_Out)
	);
	Batch_Norm bn_kernel64(
		.Data_A(32'b00111110111001011011000001101001),
		.Data_B(32'b00111111001011011001111111110010),
		.Data_In(add_k64_Data_Out),
		.Valid_In(add_kernel64_Valid_Out),
		.Data_Out(bn64_Data_Out),
		.Valid_Out(bn64_Valid_Out)
	);
	Relu_Core rl_kernel64(
		.Data_In(bn64_Data_Out),
		.Valid_In(bn64_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(rl64_Valid_Out)
	);

endmodule