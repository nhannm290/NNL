module Test_Global_AVG (
    ports
);
    
endmodule