module Depthwise_Part1_Separable_64CHANNEL_Layer6 #(
    parameter DATA_WIDHT = 32, 
    parameter IMG_WIDHT = 44,
    parameter IMG_HEIGHT =44
)
(
    input [DATA_WIDHT*64-1:0] Data_In,
    input clk,
    input rst,
    input Valid_In,
    output [DATA_WIDHT*64-1:0] Data_Out,
    output Valid_Out

);
	wire CHANNEL1_Valid_Out, CHANNEL2_Valid_Out, CHANNEL3_Valid_Out, CHANNEL4_Valid_Out, CHANNEL5_Valid_Out, CHANNEL6_Valid_Out, CHANNEL7_Valid_Out, CHANNEL8_Valid_Out, CHANNEL9_Valid_Out, CHANNEL10_Valid_Out, CHANNEL11_Valid_Out, CHANNEL12_Valid_Out, CHANNEL13_Valid_Out, CHANNEL14_Valid_Out, CHANNEL15_Valid_Out, CHANNEL16_Valid_Out, CHANNEL17_Valid_Out, CHANNEL18_Valid_Out, CHANNEL19_Valid_Out, CHANNEL20_Valid_Out, CHANNEL21_Valid_Out, CHANNEL22_Valid_Out, CHANNEL23_Valid_Out, CHANNEL24_Valid_Out,CHANNEL25_Valid_Out,CHANNEL26_Valid_Out,CHANNEL27_Valid_Out,CHANNEL28_Valid_Out,CHANNEL29_Valid_Out,CHANNEL30_Valid_Out,CHANNEL31_Valid_Out,CHANNEL32_Valid_Out,CHANNEL33_Valid_Out,CHANNEL34_Valid_Out,CHANNEL35_Valid_Out,CHANNEL36_Valid_Out,CHANNEL37_Valid_Out,CHANNEL38_Valid_Out,CHANNEL39_Valid_Out,CHANNEL40_Valid_Out,CHANNEL41_Valid_Out,CHANNEL42_Valid_Out,CHANNEL43_Valid_Out,CHANNEL44_Valid_Out,CHANNEL45_Valid_Out,CHANNEL46_Valid_Out,CHANNEL47_Valid_Out,CHANNEL48_Valid_Out,CHANNEL49_Valid_Out,CHANNEL50_Valid_Out,CHANNEL51_Valid_Out,CHANNEL52_Valid_Out,CHANNEL53_Valid_Out,CHANNEL54_Valid_Out,CHANNEL55_Valid_Out,CHANNEL56_Valid_Out,CHANNEL57_Valid_Out,CHANNEL58_Valid_Out,CHANNEL59_Valid_Out,CHANNEL60_Valid_Out,CHANNEL61_Valid_Out,CHANNEL62_Valid_Out,CHANNEL63_Valid_Out,CHANNEL64_Valid_Out;

	assign Valid_Out= CHANNEL1_Valid_Out & CHANNEL2_Valid_Out & CHANNEL3_Valid_Out & CHANNEL4_Valid_Out & CHANNEL5_Valid_Out & CHANNEL6_Valid_Out & CHANNEL7_Valid_Out & CHANNEL8_Valid_Out & CHANNEL9_Valid_Out & CHANNEL10_Valid_Out & CHANNEL11_Valid_Out & CHANNEL12_Valid_Out & CHANNEL13_Valid_Out & CHANNEL14_Valid_Out & CHANNEL15_Valid_Out & CHANNEL16_Valid_Out & CHANNEL17_Valid_Out & CHANNEL18_Valid_Out & CHANNEL19_Valid_Out & CHANNEL20_Valid_Out & CHANNEL21_Valid_Out & CHANNEL22_Valid_Out& CHANNEL23_Valid_Out& CHANNEL24_Valid_Out&CHANNEL25_Valid_Out&CHANNEL26_Valid_Out&CHANNEL27_Valid_Out&CHANNEL28_Valid_Out&CHANNEL29_Valid_Out&CHANNEL30_Valid_Out&CHANNEL31_Valid_Out&CHANNEL32_Valid_Out&CHANNEL33_Valid_Out&CHANNEL34_Valid_Out&CHANNEL35_Valid_Out&CHANNEL36_Valid_Out&CHANNEL37_Valid_Out&CHANNEL38_Valid_Out&CHANNEL39_Valid_Out&CHANNEL40_Valid_Out&CHANNEL41_Valid_Out&CHANNEL42_Valid_Out&CHANNEL43_Valid_Out&CHANNEL44_Valid_Out&CHANNEL45_Valid_Out&CHANNEL46_Valid_Out&CHANNEL47_Valid_Out&CHANNEL48_Valid_Out&CHANNEL49_Valid_Out&CHANNEL50_Valid_Out&CHANNEL51_Valid_Out&CHANNEL52_Valid_Out&CHANNEL53_Valid_Out&CHANNEL54_Valid_Out&CHANNEL55_Valid_Out&CHANNEL56_Valid_Out&CHANNEL57_Valid_Out&CHANNEL58_Valid_Out&CHANNEL59_Valid_Out&CHANNEL60_Valid_Out&CHANNEL61_Valid_Out&CHANNEL62_Valid_Out&CHANNEL63_Valid_Out&CHANNEL64_Valid_Out;

	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL1 (
			.Data_In(Data_In[DATA_WIDHT-1:0]),
			.Kernel0(32'b00111110111101111111011101111000),
			.Kernel1(32'b00111101111010001100010010001100),
			.Kernel2(32'b00111101111100101000100001111011),
			.Kernel3(32'b00111111000100101010100111110110),
			.Kernel4(32'b00111110101100010100011111000001),
			.Kernel5(32'b00111110100011101100100001000011),
			.Kernel6(32'b00111110110100011001010110001011),
			.Kernel7(32'b00111110001101000001001110010111),
			.Kernel8(32'b00111110010111010111101010000000),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT-1:0]),
			.Valid_Out(CHANNEL1_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL2 (
			.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
			.Kernel0(32'b00111110110110000001010110111001),
			.Kernel1(32'b10111101001001011011101010100110),
			.Kernel2(32'b00111101100110100111011110011111),
			.Kernel3(32'b00111110101011001111001000100010),
			.Kernel4(32'b00111101000001111111001010010110),
			.Kernel5(32'b00111110100001111011001010110110),
			.Kernel6(32'b00111110110011001000101001110100),
			.Kernel7(32'b00111111000101010100111101001001),
			.Kernel8(32'b00111111001111010100110001000111),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*2-1:DATA_WIDHT]),
			.Valid_Out(CHANNEL2_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL3 (
			.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
			.Kernel0(32'b00111111001100011111001100011100),
			.Kernel1(32'b00111100101010100001110111111001),
			.Kernel2(32'b10111101010000101110100110000001),
			.Kernel3(32'b00111110111000000010010101011010),
			.Kernel4(32'b00111110100000011001011001100010),
			.Kernel5(32'b00111110101111011111000010000011),
			.Kernel6(32'b00111110110111010010110011101010),
			.Kernel7(32'b00111110001100010100111111000101),
			.Kernel8(32'b00111100010101101011111101011000),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*3-1:DATA_WIDHT*2]),
			.Valid_Out(CHANNEL3_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL4 (
			.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
			.Kernel0(32'b10111110101011111100000110011101),
			.Kernel1(32'b10111110001101100100110000110001),
			.Kernel2(32'b10111110111011101001001010000010),
			.Kernel3(32'b10111110011111100101000101001101),
			.Kernel4(32'b10111101010011010100010011001101),
			.Kernel5(32'b10111110111111101010010101110111),
			.Kernel6(32'b10111110000001111010111001111000),
			.Kernel7(32'b10111101101010111110011000101100),
			.Kernel8(32'b00111011010011110011001011100110),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*4-1:DATA_WIDHT*3]),
			.Valid_Out(CHANNEL4_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL5 (
			.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
			.Kernel0(32'b10111100101010100001111101110000),
			.Kernel1(32'b10111101101001001101000011111101),
			.Kernel2(32'b00111110001000010001101010011110),
			.Kernel3(32'b00111110100000101101000001110010),
			.Kernel4(32'b00111110110010010000101100110110),
			.Kernel5(32'b00111101000001100111010100011011),
			.Kernel6(32'b00111111001000100010111011100100),
			.Kernel7(32'b00111111001001110110100100110000),
			.Kernel8(32'b00111111010010000000110111101011),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*5-1:DATA_WIDHT*4]),
			.Valid_Out(CHANNEL5_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL6 (
			.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
			.Kernel0(32'b00111110100111011101001100001110),
			.Kernel1(32'b00111110110100010001001111101000),
			.Kernel2(32'b00111111000011100111001111111111),
			.Kernel3(32'b10110111100100011110101101000000),
			.Kernel4(32'b10111100110010111011100000110110),
			.Kernel5(32'b10111101100001110110011000010010),
			.Kernel6(32'b10111111001111110110110000111010),
			.Kernel7(32'b10111110111010000101010110000100),
			.Kernel8(32'b10111111001110001110100011001011),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*6-1:DATA_WIDHT*5]),
			.Valid_Out(CHANNEL6_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL7 (
			.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
			.Kernel0(32'b00111111000100101001000111110010),
			.Kernel1(32'b00111110101111011010010110100110),
			.Kernel2(32'b10111101000011011011100000001010),
			.Kernel3(32'b00111101000001010010011010010011),
			.Kernel4(32'b00111110101000000010001100110110),
			.Kernel5(32'b00111110010110111010110001110011),
			.Kernel6(32'b10111101111110010100110010100011),
			.Kernel7(32'b10111101010001010001011010000101),
			.Kernel8(32'b10111111000101100101100001101011),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*7-1:DATA_WIDHT*6]),
			.Valid_Out(CHANNEL7_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL8 (
			.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
			.Kernel0(32'b10111111001001101101100110100001),
			.Kernel1(32'b10111110111011010010111110010010),
			.Kernel2(32'b10111111001100011011000010000100),
			.Kernel3(32'b10111110110110010110111110001010),
			.Kernel4(32'b00111101111110111101101101100000),
			.Kernel5(32'b10111101111010001011010000110101),
			.Kernel6(32'b00111110110111100110110011110101),
			.Kernel7(32'b00111110001011001011000001110101),
			.Kernel8(32'b00111101111001010010001101110111),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*8-1:DATA_WIDHT*7]),
			.Valid_Out(CHANNEL8_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL9 (
			.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
			.Kernel0(32'b10111110010100111100110001001100),
			.Kernel1(32'b10111101110110100010101000000001),
			.Kernel2(32'b10111110100110010100111101111000),
			.Kernel3(32'b10111110100001001110010000010010),
			.Kernel4(32'b10111101000010101101110010111000),
			.Kernel5(32'b10111101010101111101011011100001),
			.Kernel6(32'b00111111001000000110101010101000),
			.Kernel7(32'b00111110110011111010110101000110),
			.Kernel8(32'b00111111010111111100101011000100),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*9-1:DATA_WIDHT*8]),
			.Valid_Out(CHANNEL9_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL10 (
			.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
			.Kernel0(32'b10111111001101011000110000101101),
			.Kernel1(32'b10111101111100111001100010101011),
			.Kernel2(32'b10111110010011011000000101101011),
			.Kernel3(32'b10111110011111001001001101110110),
			.Kernel4(32'b00111110011101010101110011001010),
			.Kernel5(32'b10111110010111110000000001111000),
			.Kernel6(32'b00111111010001101111101111011001),
			.Kernel7(32'b00111110111010111100100001110110),
			.Kernel8(32'b00111111001010001100110001101100),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*10-1:DATA_WIDHT*9]),
			.Valid_Out(CHANNEL10_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL11 (
			.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
			.Kernel0(32'b00111101111100000001000001011111),
			.Kernel1(32'b00111111000010110110100011100111),
			.Kernel2(32'b00111110111100100110001111001001),
			.Kernel3(32'b10111110011111001010000101110000),
			.Kernel4(32'b10111110011011011100111110101001),
			.Kernel5(32'b10111110010100000101010010110110),
			.Kernel6(32'b10111110110010111101001101111100),
			.Kernel7(32'b10111110110100010011100111100111),
			.Kernel8(32'b10111110110001011101110110011010),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*11-1:DATA_WIDHT*10]),
			.Valid_Out(CHANNEL11_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL12 (
			.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
			.Kernel0(32'b10111111000000001110011010100110),
			.Kernel1(32'b10111111000101111101110001011111),
			.Kernel2(32'b10111111010101111101100000110100),
			.Kernel3(32'b00111110101001011110101011011011),
			.Kernel4(32'b00111110000100001011111001101001),
			.Kernel5(32'b10111110001101010100011101001000),
			.Kernel6(32'b00111110111001100010100111110010),
			.Kernel7(32'b00111111000111001101000100101111),
			.Kernel8(32'b00111110101111101111001111000111),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*12-1:DATA_WIDHT*11]),
			.Valid_Out(CHANNEL12_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL13 (
			.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
			.Kernel0(32'b00111111000100110010010010111100),
			.Kernel1(32'b10111101000111100101010011101110),
			.Kernel2(32'b00111110100110011110111101100100),
			.Kernel3(32'b00111110001101000111100110011111),
			.Kernel4(32'b10111011111000110000001101100011),
			.Kernel5(32'b10111101101111010011100001101101),
			.Kernel6(32'b00111111001101110001011100111111),
			.Kernel7(32'b00111110111111000000010011101011),
			.Kernel8(32'b00111110111000001111010011010110),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*13-1:DATA_WIDHT*12]),
			.Valid_Out(CHANNEL13_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL14 (
			.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
			.Kernel0(32'b10111111000101111110001111110000),
			.Kernel1(32'b10111110100010101111000011110010),
			.Kernel2(32'b00111111000001100110100011010010),
			.Kernel3(32'b10111110101101001000011100011001),
			.Kernel4(32'b00111101101011101010000100111011),
			.Kernel5(32'b00111110111000010111000010101011),
			.Kernel6(32'b00111101000000100110101000111110),
			.Kernel7(32'b00111111000010010000101110111101),
			.Kernel8(32'b00111111010000000011101001010110),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*14-1:DATA_WIDHT*13]),
			.Valid_Out(CHANNEL14_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL15 (
			.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
			.Kernel0(32'b10111110010010100010011000011111),
			.Kernel1(32'b00111110101010001001001011011100),
			.Kernel2(32'b00111100010010011001010100000111),
			.Kernel3(32'b10111110101001011000010101001111),
			.Kernel4(32'b00111101100001001001111101001011),
			.Kernel5(32'b00111110001011010000100100010111),
			.Kernel6(32'b10111111010011111101101100111011),
			.Kernel7(32'b10111111001000101010001101101101),
			.Kernel8(32'b10111110110111100000110110110101),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*15-1:DATA_WIDHT*14]),
			.Valid_Out(CHANNEL15_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL16 (
			.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
			.Kernel0(32'b00111101100010001100001001110001),
			.Kernel1(32'b00111100110100000000110011110111),
			.Kernel2(32'b00111110000001010110010111011110),
			.Kernel3(32'b00111110011001010011010000101001),
			.Kernel4(32'b00111101000101111010101001001100),
			.Kernel5(32'b00111101000010010010110000000010),
			.Kernel6(32'b00111111001000011100011101000001),
			.Kernel7(32'b00111110100001011000101001101111),
			.Kernel8(32'b00111111001101100010000100100000),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*16-1:DATA_WIDHT*15]),
			.Valid_Out(CHANNEL16_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL17 (
			.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
			.Kernel0(32'b00111111010010100010101110100101),
			.Kernel1(32'b00111111000001001110000111001110),
			.Kernel2(32'b00111111000001100001000011011011),
			.Kernel3(32'b00111110011110001000011110001100),
			.Kernel4(32'b10111110010100000110101011111110),
			.Kernel5(32'b10111110100010000100101011100101),
			.Kernel6(32'b10111101000101001011101111011101),
			.Kernel7(32'b10111110101110100110000101011101),
			.Kernel8(32'b10111110101100011111000011110110),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*17-1:DATA_WIDHT*16]),
			.Valid_Out(CHANNEL17_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL18 (
			.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
			.Kernel0(32'b00111110110011111010101000011101),
			.Kernel1(32'b00111110101101010100111000110011),
			.Kernel2(32'b00111110101001110101101100011000),
			.Kernel3(32'b00111111000000100100110101001000),
			.Kernel4(32'b00111110010000101010000000110100),
			.Kernel5(32'b00111110110100101010110101000100),
			.Kernel6(32'b00111110101110001000111110000000),
			.Kernel7(32'b00111101111110010010111111100110),
			.Kernel8(32'b00111110100010110100000001110011),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*18-1:DATA_WIDHT*17]),
			.Valid_Out(CHANNEL18_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL19 (
			.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
			.Kernel0(32'b10111110111001001001000001011011),
			.Kernel1(32'b10111110001010001100101110001011),
			.Kernel2(32'b10111110101011111111111000101110),
			.Kernel3(32'b10111110101111110011010011101111),
			.Kernel4(32'b10111110110001100100111111110100),
			.Kernel5(32'b10111110010011011110000110110001),
			.Kernel6(32'b00111111000011110000101100100101),
			.Kernel7(32'b00111110111010010010111100110000),
			.Kernel8(32'b00111111001000011110110010110111),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*19-1:DATA_WIDHT*18]),
			.Valid_Out(CHANNEL19_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL20 (
			.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
			.Kernel0(32'b10111111001011001101001101010010),
			.Kernel1(32'b10111111001000110110111101011100),
			.Kernel2(32'b10111111100000000000000100100000),
			.Kernel3(32'b00111101100010000111010110101110),
			.Kernel4(32'b00111101000101010111000011000110),
			.Kernel5(32'b10111110001001100101010010101000),
			.Kernel6(32'b00111110100001000000101101100010),
			.Kernel7(32'b00111101000011100000001001100110),
			.Kernel8(32'b10111110101011000000111111000011),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*20-1:DATA_WIDHT*19]),
			.Valid_Out(CHANNEL20_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL21 (
			.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
			.Kernel0(32'b10111110001000000101000111110101),
			.Kernel1(32'b10111110001111110001000001001100),
			.Kernel2(32'b10111110100100101000011100101100),
			.Kernel3(32'b10111110010010010110001101101111),
			.Kernel4(32'b10111110101001010011010001100101),
			.Kernel5(32'b10111110010011000100000000100000),
			.Kernel6(32'b00111111010110110010001101101110),
			.Kernel7(32'b00111110111010100100000111111110),
			.Kernel8(32'b00111111010100100010010100101000),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*21-1:DATA_WIDHT*20]),
			.Valid_Out(CHANNEL21_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL22 (
			.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
			.Kernel0(32'b10111110100101010011001101111000),
			.Kernel1(32'b10111101110001011001000010101000),
			.Kernel2(32'b10111101111000101000011000000001),
			.Kernel3(32'b10111110100100110111000001000110),
			.Kernel4(32'b00111101101111001011100001001011),
			.Kernel5(32'b10111110101000001111000011011100),
			.Kernel6(32'b10111110101111111110010001000111),
			.Kernel7(32'b10111110100111110110011110100100),
			.Kernel8(32'b10111111010000001101010100000000),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*22-1:DATA_WIDHT*21]),
			.Valid_Out(CHANNEL22_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL23 (
			.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
			.Kernel0(32'b10111111001000101111110110111111),
			.Kernel1(32'b10111111000011010010010111100001),
			.Kernel2(32'b10111111001001110111010010110101),
			.Kernel3(32'b00111110100111100111010000000111),
			.Kernel4(32'b00111110110010111101111100100011),
			.Kernel5(32'b00111110010000001010010101010001),
			.Kernel6(32'b00111110100000001111011100100011),
			.Kernel7(32'b10111100000000000100011100101101),
			.Kernel8(32'b10111101100010110111000111000001),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*23-1:DATA_WIDHT*22]),
			.Valid_Out(CHANNEL23_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL24 (
			.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
			.Kernel0(32'b00111111000000110110100110000011),
			.Kernel1(32'b10111111000001000001011111111011),
			.Kernel2(32'b10111110100111001100100101001001),
			.Kernel3(32'b00111111001101110111111101011111),
			.Kernel4(32'b00111110010000111110110111010001),
			.Kernel5(32'b10111011101001001100100001111100),
			.Kernel6(32'b00111101101000101101000111001101),
			.Kernel7(32'b10111101011010011000011011001001),
			.Kernel8(32'b10111110101110101011110100110011),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*24-1:DATA_WIDHT*23]),
			.Valid_Out(CHANNEL24_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL25 (
			.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
			.Kernel0(32'b00111110011100110000010110001110),
			.Kernel1(32'b00111110111110100100011000010110),
			.Kernel2(32'b00111110101001100111011010101111),
			.Kernel3(32'b10111110110010110110110010001100),
			.Kernel4(32'b10111110000101011011001101000010),
			.Kernel5(32'b10111101010101111011000101101010),
			.Kernel6(32'b10111111001011001110001000111100),
			.Kernel7(32'b10111110100111010110111001111101),
			.Kernel8(32'b10111110010111010011000000100110),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*25-1:DATA_WIDHT*24]),
			.Valid_Out(CHANNEL25_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL26 (
			.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
			.Kernel0(32'b10111110011100101110010110001101),
			.Kernel1(32'b00111101101101010001000100001001),
			.Kernel2(32'b00111110101011111010001101011011),
			.Kernel3(32'b00111110100111111010100010101010),
			.Kernel4(32'b00111110011010110101000100100010),
			.Kernel5(32'b00111110110011101101011110000100),
			.Kernel6(32'b00111110100010100101100111011000),
			.Kernel7(32'b00111110100111000001010001011011),
			.Kernel8(32'b00111110111101101110100101111010),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*26-1:DATA_WIDHT*25]),
			.Valid_Out(CHANNEL26_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL27 (
			.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
			.Kernel0(32'b10111110011100001001000111011001),
			.Kernel1(32'b10111110000001010110001100001010),
			.Kernel2(32'b10111110110010110111111001101110),
			.Kernel3(32'b00111110010000101010000001111000),
			.Kernel4(32'b00111110101001101111111011000000),
			.Kernel5(32'b00111111000000011101111111010110),
			.Kernel6(32'b00111110100100100111111101000101),
			.Kernel7(32'b00111110111010011100110011111101),
			.Kernel8(32'b00111111000101000000010001110100),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*27-1:DATA_WIDHT*26]),
			.Valid_Out(CHANNEL27_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL28 (
			.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
			.Kernel0(32'b00111111010000010000111110010011),
			.Kernel1(32'b00111111001000111001101101000101),
			.Kernel2(32'b00111111001110111111011000100000),
			.Kernel3(32'b00111101000000001101010011000100),
			.Kernel4(32'b00111110000011001001001100100000),
			.Kernel5(32'b00111111000001011001000011100001),
			.Kernel6(32'b10111110110101011010101101111101),
			.Kernel7(32'b00111101100011101100101110100111),
			.Kernel8(32'b00111100101001100100100011100001),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*28-1:DATA_WIDHT*27]),
			.Valid_Out(CHANNEL28_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL29 (
			.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
			.Kernel0(32'b10111110111111010000111010011110),
			.Kernel1(32'b10111110100101011010100011100011),
			.Kernel2(32'b10111111011100001011000001100101),
			.Kernel3(32'b10111101101100001001011001010000),
			.Kernel4(32'b10111110011001000011010100001110),
			.Kernel5(32'b10111110111111001001111111001000),
			.Kernel6(32'b00111110110111110110011100011111),
			.Kernel7(32'b00111110100111111100100001000110),
			.Kernel8(32'b10111101100001101101110010010000),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*29-1:DATA_WIDHT*28]),
			.Valid_Out(CHANNEL29_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL30 (
			.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
			.Kernel0(32'b00111100010001110101010010010110),
			.Kernel1(32'b10111101101110100101111001011110),
			.Kernel2(32'b00111101110011011010110101100111),
			.Kernel3(32'b00111101111000101010110010111010),
			.Kernel4(32'b00111110100001001000001000111010),
			.Kernel5(32'b10111110101011010100111101111110),
			.Kernel6(32'b00111110001110001010100011010001),
			.Kernel7(32'b10111111000011011010100001000000),
			.Kernel8(32'b10111111011110000100001111100110),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*30-1:DATA_WIDHT*29]),
			.Valid_Out(CHANNEL30_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL31 (
			.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
			.Kernel0(32'b10111110100001010011011010010001),
			.Kernel1(32'b10111100001101100111110100011001),
			.Kernel2(32'b10111110010000101101001101000101),
			.Kernel3(32'b00111110000000101001000000010101),
			.Kernel4(32'b00111110011010100101001011110110),
			.Kernel5(32'b00111110111011011010101101100100),
			.Kernel6(32'b00111111001001011001001111000000),
			.Kernel7(32'b00111110100010010100111000000001),
			.Kernel8(32'b00111111001000001010100010100111),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*31-1:DATA_WIDHT*30]),
			.Valid_Out(CHANNEL31_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL32 (
			.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
			.Kernel0(32'b10111111000111101101011100111101),
			.Kernel1(32'b10111110111110111000001010110110),
			.Kernel2(32'b10111111010001100110011011001011),
			.Kernel3(32'b00111110100101110000111100111101),
			.Kernel4(32'b10111101100101110001110010001010),
			.Kernel5(32'b00111110001110101010011111111011),
			.Kernel6(32'b00111110010100010000110110000111),
			.Kernel7(32'b00111110100100101011111010110100),
			.Kernel8(32'b00111110001110010000001110100110),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*32-1:DATA_WIDHT*31]),
			.Valid_Out(CHANNEL32_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL33 (
			.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
			.Kernel0(32'b00111101000110001101011101010011),
			.Kernel1(32'b00111100111011001000010010110010),
			.Kernel2(32'b00111101101010001100010001111001),
			.Kernel3(32'b00111110101110101010101100111011),
			.Kernel4(32'b00111101100010111010000000100101),
			.Kernel5(32'b00111110101011011111011110111011),
			.Kernel6(32'b00111111000010101111001010010000),
			.Kernel7(32'b00111110110001011111000001111111),
			.Kernel8(32'b00111111010000001010110101101110),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*33-1:DATA_WIDHT*32]),
			.Valid_Out(CHANNEL33_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL34 (
			.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
			.Kernel0(32'b00111101101010110000000110001111),
			.Kernel1(32'b10111110100011111100001011011101),
			.Kernel2(32'b10111101010000111110001010011011),
			.Kernel3(32'b10111100101010010001101011000100),
			.Kernel4(32'b10111101110111111010100101010111),
			.Kernel5(32'b00111110001110011011101100000101),
			.Kernel6(32'b00111111001011001010010101010111),
			.Kernel7(32'b00111111000001100110001011100100),
			.Kernel8(32'b00111111001000100111000010000010),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*34-1:DATA_WIDHT*33]),
			.Valid_Out(CHANNEL34_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL35 (
			.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
			.Kernel0(32'b10111110111010100010110110011101),
			.Kernel1(32'b10111110110000101111111011100100),
			.Kernel2(32'b10111111000011000010100000000011),
			.Kernel3(32'b00111101111011111110100100000110),
			.Kernel4(32'b00111110001000000011010111101000),
			.Kernel5(32'b10111101110101010101000011010011),
			.Kernel6(32'b10111110101001100111100001111100),
			.Kernel7(32'b10111110010111110001000100111000),
			.Kernel8(32'b00111100001000001001011101101000),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*35-1:DATA_WIDHT*34]),
			.Valid_Out(CHANNEL35_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL36 (
			.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
			.Kernel0(32'b00111111001011110101011010010100),
			.Kernel1(32'b00111111000001011111111111010101),
			.Kernel2(32'b00111111000100000000010011001110),
			.Kernel3(32'b10111110001011010100000100011110),
			.Kernel4(32'b10111101111010110010001011101001),
			.Kernel5(32'b10111110100000011110111011100001),
			.Kernel6(32'b10111110110011110000000110111011),
			.Kernel7(32'b10111110111101011100001010110001),
			.Kernel8(32'b10111111001001100100010010111110),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*36-1:DATA_WIDHT*35]),
			.Valid_Out(CHANNEL36_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL37 (
			.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
			.Kernel0(32'b10111110100010110110000011011000),
			.Kernel1(32'b10111110111101111110010110101101),
			.Kernel2(32'b10111110011111011111001100001011),
			.Kernel3(32'b10111110100111100100010000011011),
			.Kernel4(32'b00111110001001100101001101101101),
			.Kernel5(32'b10111110101000100000111100101110),
			.Kernel6(32'b00111110100011110101101010001001),
			.Kernel7(32'b10111110010000110110001001111110),
			.Kernel8(32'b10111110000011101100011000011000),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*37-1:DATA_WIDHT*36]),
			.Valid_Out(CHANNEL37_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL38 (
			.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
			.Kernel0(32'b00111110110011001001010000110111),
			.Kernel1(32'b00111110000101011110010001000100),
			.Kernel2(32'b10111101110011011100011101010111),
			.Kernel3(32'b00111111001100101100001100100111),
			.Kernel4(32'b10111110011000000011010001000001),
			.Kernel5(32'b10111111001100111100100100000110),
			.Kernel6(32'b00111111001101011100001101000001),
			.Kernel7(32'b10111110000101010011101111100110),
			.Kernel8(32'b10111111000100011111110001000101),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*38-1:DATA_WIDHT*37]),
			.Valid_Out(CHANNEL38_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL39 (
			.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
			.Kernel0(32'b10111110110000100011111010110000),
			.Kernel1(32'b10111110011011000010010000101000),
			.Kernel2(32'b10111110000011100101100101001000),
			.Kernel3(32'b10111110100001100110001011001000),
			.Kernel4(32'b10111101110100111000101100101001),
			.Kernel5(32'b10111101110110111101101001100011),
			.Kernel6(32'b10111110110101111100000011001011),
			.Kernel7(32'b00111110001101000010100110100101),
			.Kernel8(32'b10111100111110011111110001001110),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*39-1:DATA_WIDHT*38]),
			.Valid_Out(CHANNEL39_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL40 (
			.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
			.Kernel0(32'b00111110000010110010101010001101),
			.Kernel1(32'b00111011000010011001011000110110),
			.Kernel2(32'b00111110000011101111011000010000),
			.Kernel3(32'b00111110100101001110001001101101),
			.Kernel4(32'b10111101010010110010010101100100),
			.Kernel5(32'b00111110010001101001100010101001),
			.Kernel6(32'b00111111000101100011101001110010),
			.Kernel7(32'b00111110101010010010100011010010),
			.Kernel8(32'b00111111001110111011111111101101),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*40-1:DATA_WIDHT*39]),
			.Valid_Out(CHANNEL40_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL41 (
			.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
			.Kernel0(32'b00111100111001010101111111101110),
			.Kernel1(32'b10111110101111111001000101110001),
			.Kernel2(32'b10111111000101111011110110101111),
			.Kernel3(32'b00111101101010100000111010010101),
			.Kernel4(32'b00111110100010100110010001001000),
			.Kernel5(32'b10111101100100000011100000101100),
			.Kernel6(32'b10111110100111000010110100001001),
			.Kernel7(32'b00111100000011110100001010100001),
			.Kernel8(32'b10111110101111010011100111001101),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*41-1:DATA_WIDHT*40]),
			.Valid_Out(CHANNEL41_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL42 (
			.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
			.Kernel0(32'b00111110110001110110011000000010),
			.Kernel1(32'b00111111000101100001111110111110),
			.Kernel2(32'b00111111000110101010100010101111),
			.Kernel3(32'b10111110100000101011101011001000),
			.Kernel4(32'b00111101101011011111100111100000),
			.Kernel5(32'b00111110010010001001101111000100),
			.Kernel6(32'b00111110101010100110010111001000),
			.Kernel7(32'b00111110011110111011101110001100),
			.Kernel8(32'b00111110001000000101100010001011),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*42-1:DATA_WIDHT*41]),
			.Valid_Out(CHANNEL42_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL43 (
			.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
			.Kernel0(32'b10111111011011010010101011001000),
			.Kernel1(32'b10111110111111010010111101000011),
			.Kernel2(32'b10111110100100111110111101100010),
			.Kernel3(32'b00111101110001111010000101010101),
			.Kernel4(32'b10111110010010011101111001011110),
			.Kernel5(32'b10111110100110101010110110010001),
			.Kernel6(32'b00111111000001100010100001100001),
			.Kernel7(32'b00111111000101110110010111000011),
			.Kernel8(32'b00111111000100011000111111101110),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*43-1:DATA_WIDHT*42]),
			.Valid_Out(CHANNEL43_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL44 (
			.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
			.Kernel0(32'b00111111011000111100110011110011),
			.Kernel1(32'b00111110110101010101001011110111),
			.Kernel2(32'b00111111001111011101011010001111),
			.Kernel3(32'b10111101100100110001000111011011),
			.Kernel4(32'b00111101100110111101100111011011),
			.Kernel5(32'b10111101111111001111101101110010),
			.Kernel6(32'b10111110111101101001011111001111),
			.Kernel7(32'b10111111000111100010001000101101),
			.Kernel8(32'b10111110100000001100100001111010),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*44-1:DATA_WIDHT*43]),
			.Valid_Out(CHANNEL44_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL45 (
			.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
			.Kernel0(32'b10111111000101101010111010100101),
			.Kernel1(32'b10111110111011011111001111110010),
			.Kernel2(32'b10111110001011100101000101010110),
			.Kernel3(32'b10111110011101010100000100111110),
			.Kernel4(32'b10111110011101001111011001011101),
			.Kernel5(32'b10111110001100110001110001111000),
			.Kernel6(32'b10111101000111010111010001000111),
			.Kernel7(32'b10111101110001111100101011010000),
			.Kernel8(32'b10111101110000100101100000011111),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*45-1:DATA_WIDHT*44]),
			.Valid_Out(CHANNEL45_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL46 (
			.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
			.Kernel0(32'b10111111000100000010010100010110),
			.Kernel1(32'b10111111000101010100000101011011),
			.Kernel2(32'b10111111010111011011110000100111),
			.Kernel3(32'b00111101111000111111011110100010),
			.Kernel4(32'b00111101100111001101010000000101),
			.Kernel5(32'b10111110100001100001111101111110),
			.Kernel6(32'b00111110101111011001000111011001),
			.Kernel7(32'b00111110101001111000000100000100),
			.Kernel8(32'b10111101110010000000011000101010),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*46-1:DATA_WIDHT*45]),
			.Valid_Out(CHANNEL46_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL47 (
			.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
			.Kernel0(32'b00111111011000011100001000111111),
			.Kernel1(32'b00111111000010011100001010100101),
			.Kernel2(32'b00111110100111000010101000111101),
			.Kernel3(32'b00111110111110100000010110110000),
			.Kernel4(32'b10111100010011110010001110000010),
			.Kernel5(32'b00111110001110101000111000000010),
			.Kernel6(32'b10111110001011000001011011100011),
			.Kernel7(32'b10111110001010100111111110110110),
			.Kernel8(32'b00111101101111000001000101101011),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*47-1:DATA_WIDHT*46]),
			.Valid_Out(CHANNEL47_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL48 (
			.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
			.Kernel0(32'b00111111011000111011110011100001),
			.Kernel1(32'b00111111001001101110100110100010),
			.Kernel2(32'b00111111010011110111111111101101),
			.Kernel3(32'b10111110010100001010110001001111),
			.Kernel4(32'b10111110011011001010110100010011),
			.Kernel5(32'b00111101101110100001001110110111),
			.Kernel6(32'b10111101010111000110100010010010),
			.Kernel7(32'b10111110100000001010010011000110),
			.Kernel8(32'b10111110100111001100000100101111),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*48-1:DATA_WIDHT*47]),
			.Valid_Out(CHANNEL48_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL49 (
			.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
			.Kernel0(32'b00111110111100010001001000100001),
			.Kernel1(32'b00111110110101000010111011100010),
			.Kernel2(32'b00111111001100000111100000111000),
			.Kernel3(32'b00111110010100101100011100000100),
			.Kernel4(32'b00111101111111011101011000111100),
			.Kernel5(32'b00111101100011101110110100010001),
			.Kernel6(32'b10111110110010010001011111101000),
			.Kernel7(32'b10111111000101010111010000100101),
			.Kernel8(32'b10111111001110001000110000001011),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*49-1:DATA_WIDHT*48]),
			.Valid_Out(CHANNEL49_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL50 (
			.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
			.Kernel0(32'b00111111001010101010001110001001),
			.Kernel1(32'b00111110110111111100111110101111),
			.Kernel2(32'b00111111001100110010101000110000),
			.Kernel3(32'b00111110011010110000100001010100),
			.Kernel4(32'b00111110010111100111011001001011),
			.Kernel5(32'b00111110100111000110000000111000),
			.Kernel6(32'b00111110000111001111111000001110),
			.Kernel7(32'b10111110101111100111010000010000),
			.Kernel8(32'b00111101110101101110111010111111),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*50-1:DATA_WIDHT*49]),
			.Valid_Out(CHANNEL50_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL51 (
			.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
			.Kernel0(32'b10111110010101110000010101101001),
			.Kernel1(32'b00111101101101011010101000011101),
			.Kernel2(32'b00111100111011011010100011110111),
			.Kernel3(32'b10111101111110100101111011100001),
			.Kernel4(32'b00111101001001101101100000000100),
			.Kernel5(32'b00111101000100101011000110101010),
			.Kernel6(32'b10111111010011100001101011000111),
			.Kernel7(32'b10111111001100011101011001001111),
			.Kernel8(32'b10111111001110100100101111000101),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*51-1:DATA_WIDHT*50]),
			.Valid_Out(CHANNEL51_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL52 (
			.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
			.Kernel0(32'b00111111001101001010010011110000),
			.Kernel1(32'b00111111000001000001101001110111),
			.Kernel2(32'b00111111100010000101100110000010),
			.Kernel3(32'b10111110000010001011111101100000),
			.Kernel4(32'b00111100010000000110111000100001),
			.Kernel5(32'b00111110001001001100111000111100),
			.Kernel6(32'b10111101001100111101111111010110),
			.Kernel7(32'b10111110011011001111100110111000),
			.Kernel8(32'b00111110110111010100101000001110),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*52-1:DATA_WIDHT*51]),
			.Valid_Out(CHANNEL52_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL53 (
			.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
			.Kernel0(32'b00111111010110100111010110100111),
			.Kernel1(32'b00111111000101000000110000000000),
			.Kernel2(32'b00111110111101010111101000000000),
			.Kernel3(32'b00111110111000011001010100111100),
			.Kernel4(32'b10111101110100010111000011001101),
			.Kernel5(32'b10111101111001110001001101100110),
			.Kernel6(32'b10111101111000001101111011111001),
			.Kernel7(32'b10111110111001101001010011011000),
			.Kernel8(32'b10111110011100001010010001011011),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*53-1:DATA_WIDHT*52]),
			.Valid_Out(CHANNEL53_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL54 (
			.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
			.Kernel0(32'b00111110001100110110110001101011),
			.Kernel1(32'b00111101111111110101010111010010),
			.Kernel2(32'b10111110000101010101000110001101),
			.Kernel3(32'b00111101110100100000110110111010),
			.Kernel4(32'b10111110011000001100011011011000),
			.Kernel5(32'b00111101010111011101010100111100),
			.Kernel6(32'b10111111000101101000001001001010),
			.Kernel7(32'b10111110111011100111100101101011),
			.Kernel8(32'b10111111000011111100011000100110),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*54-1:DATA_WIDHT*53]),
			.Valid_Out(CHANNEL54_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL55 (
			.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
			.Kernel0(32'b00111111001000111111011010000111),
			.Kernel1(32'b00111110101111000111101001000000),
			.Kernel2(32'b00111111000101100001011011100111),
			.Kernel3(32'b00111110100100100100000000001101),
			.Kernel4(32'b00111110100100010110101111111100),
			.Kernel5(32'b00111101010011100000001110110101),
			.Kernel6(32'b00111110100010001111010101010000),
			.Kernel7(32'b00111110011111111010010011110000),
			.Kernel8(32'b00111101101011101010001010010110),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*55-1:DATA_WIDHT*54]),
			.Valid_Out(CHANNEL55_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL56 (
			.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
			.Kernel0(32'b00111110101000000010111110111001),
			.Kernel1(32'b00111110110001111010010111010001),
			.Kernel2(32'b00111110111110011110101001100011),
			.Kernel3(32'b10111101101111110000100001010100),
			.Kernel4(32'b10111101111011100101110101010001),
			.Kernel5(32'b00111101010111101110111111010100),
			.Kernel6(32'b10111111011001101000101010111100),
			.Kernel7(32'b10111110100010011100001010110010),
			.Kernel8(32'b10111111001000101000011011101001),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*56-1:DATA_WIDHT*55]),
			.Valid_Out(CHANNEL56_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL57 (
			.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
			.Kernel0(32'b10111111010000001110111110101011),
			.Kernel1(32'b10111110001001101101101000001010),
			.Kernel2(32'b10111111010000111000001111001111),
			.Kernel3(32'b10111101101111000110000100100101),
			.Kernel4(32'b10111110100001010001101011110010),
			.Kernel5(32'b00111101011000010111100011011000),
			.Kernel6(32'b00111100001000001100101011010101),
			.Kernel7(32'b10111101011000110011110011010010),
			.Kernel8(32'b00111101001000000000001011100101),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*57-1:DATA_WIDHT*56]),
			.Valid_Out(CHANNEL57_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL58 (
			.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
			.Kernel0(32'b10111110011100101111111110110010),
			.Kernel1(32'b10111101010111101001101100111100),
			.Kernel2(32'b10111110011001010011100001011110),
			.Kernel3(32'b00111101010011011001011000110000),
			.Kernel4(32'b10111100101001100110011101100100),
			.Kernel5(32'b10111110001101101000010101100011),
			.Kernel6(32'b10111111000110010001001110001100),
			.Kernel7(32'b10111111000101111110111010101101),
			.Kernel8(32'b10111111001110000001011010111110),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*58-1:DATA_WIDHT*57]),
			.Valid_Out(CHANNEL58_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL59 (
			.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
			.Kernel0(32'b10111110100001111111101101100110),
			.Kernel1(32'b10111110101010000100001011001111),
			.Kernel2(32'b10111111001010001010011111011101),
			.Kernel3(32'b00111111010000011000011010011101),
			.Kernel4(32'b00111111000010010111110101001100),
			.Kernel5(32'b00111110111101111011010001000001),
			.Kernel6(32'b00111110110111101111101000011111),
			.Kernel7(32'b00111110101100010101111010001000),
			.Kernel8(32'b00111110100010111000100001101111),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*59-1:DATA_WIDHT*58]),
			.Valid_Out(CHANNEL59_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL60 (
			.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
			.Kernel0(32'b00111110111000101001100110011000),
			.Kernel1(32'b00111111000010000011010110100100),
			.Kernel2(32'b00111110111110111100100111100011),
			.Kernel3(32'b10111101111101100110101100000011),
			.Kernel4(32'b10111110011000100111110010010101),
			.Kernel5(32'b00111111000011001111000001000010),
			.Kernel6(32'b10111110110111111101001010101011),
			.Kernel7(32'b10111110101101011111011111110010),
			.Kernel8(32'b00111100100001000110001101011001),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*60-1:DATA_WIDHT*59]),
			.Valid_Out(CHANNEL60_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL61 (
			.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
			.Kernel0(32'b10111100001011100101101000001110),
			.Kernel1(32'b00111101111000100001101011000100),
			.Kernel2(32'b00111100000111100101101100111100),
			.Kernel3(32'b00111110111011111010010111100000),
			.Kernel4(32'b10111101101111011001010010111101),
			.Kernel5(32'b00111110100010001011000011111101),
			.Kernel6(32'b00111111010011111110010100110011),
			.Kernel7(32'b00111110111101100111101010111011),
			.Kernel8(32'b00111111011111100000111010011001),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*61-1:DATA_WIDHT*60]),
			.Valid_Out(CHANNEL61_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL62 (
			.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
			.Kernel0(32'b00111111001001011010100001101000),
			.Kernel1(32'b00111110010001110001100100111000),
			.Kernel2(32'b00111111001011111100100000011010),
			.Kernel3(32'b00111101101111010110110100111011),
			.Kernel4(32'b00111101111000110101111000011110),
			.Kernel5(32'b00111110011101011100100101001001),
			.Kernel6(32'b00111110001010011100100010110101),
			.Kernel7(32'b00111110101101100010101111100010),
			.Kernel8(32'b00111110011100011000010010111010),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*62-1:DATA_WIDHT*61]),
			.Valid_Out(CHANNEL62_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL63 (
			.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
			.Kernel0(32'b10111111000010000111000011010100),
			.Kernel1(32'b10111110001010111001111010101101),
			.Kernel2(32'b10111110111101100000110001000011),
			.Kernel3(32'b10111110011000001100110010101110),
			.Kernel4(32'b10111110001010111100110011111110),
			.Kernel5(32'b10111110001110101010001101111010),
			.Kernel6(32'b10111110000100100001110110001011),
			.Kernel7(32'b10111110100100101100000101011111),
			.Kernel8(32'b10111110101110000110011001010001),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*63-1:DATA_WIDHT*62]),
			.Valid_Out(CHANNEL63_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL64 (
			.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
			.Kernel0(32'b00111110001010001000101001000001),
			.Kernel1(32'b10111110101100100101101111000100),
			.Kernel2(32'b10111110111001111000011110111100),
			.Kernel3(32'b00111111000100011011001100100001),
			.Kernel4(32'b10111110000000101111101010010000),
			.Kernel5(32'b10111100010011101111111010111010),
			.Kernel6(32'b00111111000101111111011011010000),
			.Kernel7(32'b00111110110010011110001111001011),
			.Kernel8(32'b00111110100011100000101110010100),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*64-1:DATA_WIDHT*63]),
			.Valid_Out(CHANNEL64_Valid_Out)
		);

    
endmodule