module Depthwise_Part1_Separable_128CHANNEL_Layer6 #(
    parameter DATA_WIDHT = 32, 
    parameter IMG_WIDHT = 44,
    parameter IMG_HEIGHT =44
)
(
    input [DATA_WIDHT*128-1:0] Data_In,
    input clk,
    input rst,
    input Valid_In,
    output [DATA_WIDHT*128-1:0] Data_Out,
    output Valid_Out

);
	wire CHANNEL1_Valid_Out, CHANNEL2_Valid_Out, CHANNEL3_Valid_Out, CHANNEL4_Valid_Out, CHANNEL5_Valid_Out, CHANNEL6_Valid_Out, CHANNEL7_Valid_Out, CHANNEL8_Valid_Out, CHANNEL9_Valid_Out, CHANNEL10_Valid_Out, CHANNEL11_Valid_Out, CHANNEL12_Valid_Out, CHANNEL13_Valid_Out, CHANNEL14_Valid_Out, CHANNEL15_Valid_Out, CHANNEL16_Valid_Out, CHANNEL17_Valid_Out, CHANNEL18_Valid_Out, CHANNEL19_Valid_Out, CHANNEL20_Valid_Out, CHANNEL21_Valid_Out, CHANNEL22_Valid_Out, CHANNEL23_Valid_Out, CHANNEL24_Valid_Out, CHANNEL25_Valid_Out, CHANNEL26_Valid_Out, CHANNEL27_Valid_Out, CHANNEL28_Valid_Out, CHANNEL29_Valid_Out, CHANNEL30_Valid_Out, CHANNEL31_Valid_Out, CHANNEL32_Valid_Out, CHANNEL33_Valid_Out, CHANNEL34_Valid_Out, CHANNEL35_Valid_Out, CHANNEL36_Valid_Out, CHANNEL37_Valid_Out, CHANNEL38_Valid_Out, CHANNEL39_Valid_Out, CHANNEL40_Valid_Out, CHANNEL41_Valid_Out, CHANNEL42_Valid_Out, CHANNEL43_Valid_Out, CHANNEL44_Valid_Out, CHANNEL45_Valid_Out, CHANNEL46_Valid_Out, CHANNEL47_Valid_Out, CHANNEL48_Valid_Out, CHANNEL49_Valid_Out, CHANNEL50_Valid_Out, CHANNEL51_Valid_Out, CHANNEL52_Valid_Out, CHANNEL53_Valid_Out, CHANNEL54_Valid_Out, CHANNEL55_Valid_Out, CHANNEL56_Valid_Out, CHANNEL57_Valid_Out, CHANNEL58_Valid_Out, CHANNEL59_Valid_Out, CHANNEL60_Valid_Out, CHANNEL61_Valid_Out, CHANNEL62_Valid_Out, CHANNEL63_Valid_Out, CHANNEL64_Valid_Out, CHANNEL65_Valid_Out, CHANNEL66_Valid_Out, CHANNEL67_Valid_Out, CHANNEL68_Valid_Out, CHANNEL69_Valid_Out, CHANNEL70_Valid_Out, CHANNEL71_Valid_Out, CHANNEL72_Valid_Out, CHANNEL73_Valid_Out, CHANNEL74_Valid_Out, CHANNEL75_Valid_Out, CHANNEL76_Valid_Out, CHANNEL77_Valid_Out, CHANNEL78_Valid_Out, CHANNEL79_Valid_Out, CHANNEL80_Valid_Out, CHANNEL81_Valid_Out, CHANNEL82_Valid_Out, CHANNEL83_Valid_Out, CHANNEL84_Valid_Out, CHANNEL85_Valid_Out, CHANNEL86_Valid_Out, CHANNEL87_Valid_Out, CHANNEL88_Valid_Out, CHANNEL89_Valid_Out, CHANNEL90_Valid_Out, CHANNEL91_Valid_Out, CHANNEL92_Valid_Out, CHANNEL93_Valid_Out, CHANNEL94_Valid_Out, CHANNEL95_Valid_Out, CHANNEL96_Valid_Out, CHANNEL97_Valid_Out, CHANNEL98_Valid_Out, CHANNEL99_Valid_Out, CHANNEL100_Valid_Out, CHANNEL101_Valid_Out, CHANNEL102_Valid_Out, CHANNEL103_Valid_Out, CHANNEL104_Valid_Out, CHANNEL105_Valid_Out, CHANNEL106_Valid_Out, CHANNEL107_Valid_Out, CHANNEL108_Valid_Out, CHANNEL109_Valid_Out, CHANNEL110_Valid_Out, CHANNEL111_Valid_Out, CHANNEL112_Valid_Out, CHANNEL113_Valid_Out, CHANNEL114_Valid_Out, CHANNEL115_Valid_Out, CHANNEL116_Valid_Out, CHANNEL117_Valid_Out, CHANNEL118_Valid_Out, CHANNEL119_Valid_Out, CHANNEL120_Valid_Out, CHANNEL121_Valid_Out, CHANNEL122_Valid_Out, CHANNEL123_Valid_Out, CHANNEL124_Valid_Out, CHANNEL125_Valid_Out, CHANNEL126_Valid_Out, CHANNEL127_Valid_Out, CHANNEL128_Valid_Out;

	assign Valid_Out= CHANNEL1_Valid_Out & CHANNEL2_Valid_Out & CHANNEL3_Valid_Out & CHANNEL4_Valid_Out & CHANNEL5_Valid_Out & CHANNEL6_Valid_Out & CHANNEL7_Valid_Out & CHANNEL8_Valid_Out & CHANNEL9_Valid_Out & CHANNEL10_Valid_Out & CHANNEL11_Valid_Out & CHANNEL12_Valid_Out & CHANNEL13_Valid_Out & CHANNEL14_Valid_Out & CHANNEL15_Valid_Out & CHANNEL16_Valid_Out & CHANNEL17_Valid_Out & CHANNEL18_Valid_Out & CHANNEL19_Valid_Out & CHANNEL20_Valid_Out & CHANNEL21_Valid_Out & CHANNEL22_Valid_Out & CHANNEL23_Valid_Out & CHANNEL24_Valid_Out & CHANNEL25_Valid_Out & CHANNEL26_Valid_Out & CHANNEL27_Valid_Out & CHANNEL28_Valid_Out & CHANNEL29_Valid_Out & CHANNEL30_Valid_Out & CHANNEL31_Valid_Out & CHANNEL32_Valid_Out & CHANNEL33_Valid_Out & CHANNEL34_Valid_Out & CHANNEL35_Valid_Out & CHANNEL36_Valid_Out & CHANNEL37_Valid_Out & CHANNEL38_Valid_Out & CHANNEL39_Valid_Out & CHANNEL40_Valid_Out & CHANNEL41_Valid_Out & CHANNEL42_Valid_Out & CHANNEL43_Valid_Out & CHANNEL44_Valid_Out & CHANNEL45_Valid_Out & CHANNEL46_Valid_Out & CHANNEL47_Valid_Out & CHANNEL48_Valid_Out & CHANNEL49_Valid_Out & CHANNEL50_Valid_Out & CHANNEL51_Valid_Out & CHANNEL52_Valid_Out & CHANNEL53_Valid_Out & CHANNEL54_Valid_Out & CHANNEL55_Valid_Out & CHANNEL56_Valid_Out & CHANNEL57_Valid_Out & CHANNEL58_Valid_Out & CHANNEL59_Valid_Out & CHANNEL60_Valid_Out & CHANNEL61_Valid_Out & CHANNEL62_Valid_Out & CHANNEL63_Valid_Out & CHANNEL64_Valid_Out & CHANNEL65_Valid_Out & CHANNEL66_Valid_Out & CHANNEL67_Valid_Out & CHANNEL68_Valid_Out & CHANNEL69_Valid_Out & CHANNEL70_Valid_Out & CHANNEL71_Valid_Out & CHANNEL72_Valid_Out & CHANNEL73_Valid_Out & CHANNEL74_Valid_Out & CHANNEL75_Valid_Out & CHANNEL76_Valid_Out & CHANNEL77_Valid_Out & CHANNEL78_Valid_Out & CHANNEL79_Valid_Out & CHANNEL80_Valid_Out & CHANNEL81_Valid_Out & CHANNEL82_Valid_Out & CHANNEL83_Valid_Out & CHANNEL84_Valid_Out & CHANNEL85_Valid_Out & CHANNEL86_Valid_Out & CHANNEL87_Valid_Out & CHANNEL88_Valid_Out & CHANNEL89_Valid_Out & CHANNEL90_Valid_Out & CHANNEL91_Valid_Out & CHANNEL92_Valid_Out & CHANNEL93_Valid_Out & CHANNEL94_Valid_Out & CHANNEL95_Valid_Out & CHANNEL96_Valid_Out & CHANNEL97_Valid_Out & CHANNEL98_Valid_Out & CHANNEL99_Valid_Out & CHANNEL100_Valid_Out & CHANNEL101_Valid_Out & CHANNEL102_Valid_Out & CHANNEL103_Valid_Out & CHANNEL104_Valid_Out & CHANNEL105_Valid_Out & CHANNEL106_Valid_Out & CHANNEL107_Valid_Out & CHANNEL108_Valid_Out & CHANNEL109_Valid_Out & CHANNEL110_Valid_Out & CHANNEL111_Valid_Out & CHANNEL112_Valid_Out & CHANNEL113_Valid_Out & CHANNEL114_Valid_Out & CHANNEL115_Valid_Out & CHANNEL116_Valid_Out & CHANNEL117_Valid_Out & CHANNEL118_Valid_Out & CHANNEL119_Valid_Out & CHANNEL120_Valid_Out & CHANNEL121_Valid_Out & CHANNEL122_Valid_Out & CHANNEL123_Valid_Out & CHANNEL124_Valid_Out & CHANNEL125_Valid_Out & CHANNEL126_Valid_Out & CHANNEL127_Valid_Out & CHANNEL128_Valid_Out;


	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL1 (
			.Data_In(Data_In[DATA_WIDHT-1:0]),
			.Kernel0(32'b10111110111011100011100010000010),
			.Kernel1(32'b10111110100011110001000100000100),
			.Kernel2(32'b10111110010011011101011000100000),
			.Kernel3(32'b10111101111110100011011110100111),
			.Kernel4(32'b10111111000000110101000110001000),
			.Kernel5(32'b10111110001110110110011011101100),
			.Kernel6(32'b10111110000111100101011101000010),
			.Kernel7(32'b10111110111011111100111100101110),
			.Kernel8(32'b10111110100100111011101000000111),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT-1:0]),
			.Valid_Out(CHANNEL1_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL2 (
			.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
			.Kernel0(32'b00111111000101000111100110001111),
			.Kernel1(32'b00111111000101100011101000001001),
			.Kernel2(32'b00111110000100111011000001100100),
			.Kernel3(32'b00111110100110110100100110111011),
			.Kernel4(32'b00111110101011000100100101001000),
			.Kernel5(32'b10111100110011010100111010011000),
			.Kernel6(32'b00111101111011010010111010011000),
			.Kernel7(32'b00111111000000000000111010000011),
			.Kernel8(32'b00111101110010111010011101010011),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*2-1:DATA_WIDHT]),
			.Valid_Out(CHANNEL2_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL3 (
			.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
			.Kernel0(32'b10111111001111111110110011010001),
			.Kernel1(32'b10111110100110111001010101101110),
			.Kernel2(32'b10111110110011111101000110001010),
			.Kernel3(32'b00111100101110100000000110001011),
			.Kernel4(32'b00111101010011011100111100101100),
			.Kernel5(32'b00111101010100001111101101001010),
			.Kernel6(32'b00111111000011110100010011000101),
			.Kernel7(32'b00111111000011011010001001101100),
			.Kernel8(32'b00111111000100001010110010101011),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*3-1:DATA_WIDHT*2]),
			.Valid_Out(CHANNEL3_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL4 (
			.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
			.Kernel0(32'b00111110111010001010001100010000),
			.Kernel1(32'b00111010111010111110001110101001),
			.Kernel2(32'b00111111001101000001111110111100),
			.Kernel3(32'b00111101010011100111101100000000),
			.Kernel4(32'b00111110100100001110111100000010),
			.Kernel5(32'b10111110001011100101010011000010),
			.Kernel6(32'b00111110011010010001110010101100),
			.Kernel7(32'b10111110011001001100110101111000),
			.Kernel8(32'b00111110001001101100111111000011),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*4-1:DATA_WIDHT*3]),
			.Valid_Out(CHANNEL4_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL5 (
			.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
			.Kernel0(32'b00111110111101010011110100001000),
			.Kernel1(32'b10111101110001100011111011111100),
			.Kernel2(32'b00111110101001111111000001100111),
			.Kernel3(32'b00111110111100001000110100110001),
			.Kernel4(32'b00111110110000010001111011101110),
			.Kernel5(32'b00111111000100000111000101111011),
			.Kernel6(32'b00111110000010010011111100110000),
			.Kernel7(32'b00111110101111101111011011001000),
			.Kernel8(32'b00111110101011001001111010101110),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*5-1:DATA_WIDHT*4]),
			.Valid_Out(CHANNEL5_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL6 (
			.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
			.Kernel0(32'b10111110111011001101100001101001),
			.Kernel1(32'b10111110100000010110001101110100),
			.Kernel2(32'b10111110111010101111010000100110),
			.Kernel3(32'b10111110100011111000110100011111),
			.Kernel4(32'b10111110111100111100010011010011),
			.Kernel5(32'b10111110101000000011101011000100),
			.Kernel6(32'b10111110011011000001000111111101),
			.Kernel7(32'b10111101101000111011100110101100),
			.Kernel8(32'b00111110000001101000100001000000),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*6-1:DATA_WIDHT*5]),
			.Valid_Out(CHANNEL6_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL7 (
			.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
			.Kernel0(32'b10111110110101110101111011100010),
			.Kernel1(32'b10111110110011010001110001110110),
			.Kernel2(32'b00111111001101010111100101010000),
			.Kernel3(32'b10111110011010001001110001110010),
			.Kernel4(32'b10111110110110100110000111001100),
			.Kernel5(32'b00111110111110110011111100011111),
			.Kernel6(32'b00111101111010010001001110100101),
			.Kernel7(32'b10111110101101010010101010101010),
			.Kernel8(32'b00111110101000111011010110101111),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*7-1:DATA_WIDHT*6]),
			.Valid_Out(CHANNEL7_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL8 (
			.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
			.Kernel0(32'b10111111000011001001011100001001),
			.Kernel1(32'b10111111000111011110010111000101),
			.Kernel2(32'b10111110111100101000001010010010),
			.Kernel3(32'b10111110110101000101000111111001),
			.Kernel4(32'b10111111000110110100010000001011),
			.Kernel5(32'b10111110001111100110100100110101),
			.Kernel6(32'b10111110100000001000000001001010),
			.Kernel7(32'b00111110010100110100001011100100),
			.Kernel8(32'b00111110011010010111101001000110),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*8-1:DATA_WIDHT*7]),
			.Valid_Out(CHANNEL8_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL9 (
			.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
			.Kernel0(32'b00111111000111010000111011011110),
			.Kernel1(32'b00111110010110101000001001111010),
			.Kernel2(32'b00111110111001000111001000011110),
			.Kernel3(32'b10111110010100111001110000111000),
			.Kernel4(32'b10111110110110101000011000000111),
			.Kernel5(32'b10111110110011110011000101110111),
			.Kernel6(32'b00111101001111111001001010011001),
			.Kernel7(32'b10111110101100111100110000111010),
			.Kernel8(32'b10111110100000111010001100000011),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*9-1:DATA_WIDHT*8]),
			.Valid_Out(CHANNEL9_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL10 (
			.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
			.Kernel0(32'b10111110101000110111111011111011),
			.Kernel1(32'b10111110100010011011110001110000),
			.Kernel2(32'b10111110101110001101111011111110),
			.Kernel3(32'b10111110101001101111011111000111),
			.Kernel4(32'b10111110100010001101110011100101),
			.Kernel5(32'b10111110101100001110100000100110),
			.Kernel6(32'b10111110101100000101111011011101),
			.Kernel7(32'b10111110011001101000100100111010),
			.Kernel8(32'b10111110101101111011100001010110),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*10-1:DATA_WIDHT*9]),
			.Valid_Out(CHANNEL10_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL11 (
			.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
			.Kernel0(32'b10111111000111001111011110110011),
			.Kernel1(32'b10111111000001010110100000001111),
			.Kernel2(32'b10111111010000101101010011011011),
			.Kernel3(32'b10111110011101101101011000110101),
			.Kernel4(32'b10111110000010100111101111000111),
			.Kernel5(32'b10111101111001000110010010110000),
			.Kernel6(32'b10111110011110111000010001011011),
			.Kernel7(32'b10111110010110101101100001001000),
			.Kernel8(32'b00111101011001111111000011100001),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*11-1:DATA_WIDHT*10]),
			.Valid_Out(CHANNEL11_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL12 (
			.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
			.Kernel0(32'b00111111000101010010010011100110),
			.Kernel1(32'b00111100111011101101010000100000),
			.Kernel2(32'b00111110001100000000101101010000),
			.Kernel3(32'b00111110100011000100001000000000),
			.Kernel4(32'b00111110110101001011011110111111),
			.Kernel5(32'b00111111000000111011101111000011),
			.Kernel6(32'b00111111001111000111001101010111),
			.Kernel7(32'b00111110100000101111001010001101),
			.Kernel8(32'b00111111001010101000011111000101),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*12-1:DATA_WIDHT*11]),
			.Valid_Out(CHANNEL12_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL13 (
			.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
			.Kernel0(32'b00111111000001001110001101101111),
			.Kernel1(32'b00111111000101000000001100111010),
			.Kernel2(32'b00111111011000000001000011001100),
			.Kernel3(32'b10111100110110110111010000111000),
			.Kernel4(32'b10111110100110010000011000101100),
			.Kernel5(32'b10111101001111100111011001011101),
			.Kernel6(32'b10111111010100100000000001110000),
			.Kernel7(32'b10111111000001011001011001111011),
			.Kernel8(32'b10111111010000011100101001011000),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*13-1:DATA_WIDHT*12]),
			.Valid_Out(CHANNEL13_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL14 (
			.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
			.Kernel0(32'b00111111001100100001011011010010),
			.Kernel1(32'b00111110011100110001011001100010),
			.Kernel2(32'b00111110111000100110010010101011),
			.Kernel3(32'b10111110101101101101110100111000),
			.Kernel4(32'b10111110001100011110110000000000),
			.Kernel5(32'b10111111000000010011001001010111),
			.Kernel6(32'b10111111010000110001101100111101),
			.Kernel7(32'b10111111000010100001100001101101),
			.Kernel8(32'b10111110011000010001001000101110),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*14-1:DATA_WIDHT*13]),
			.Valid_Out(CHANNEL14_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL15 (
			.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
			.Kernel0(32'b00111111010100110000010101110111),
			.Kernel1(32'b00111111000101111100101011100000),
			.Kernel2(32'b00111111010010000010001111111001),
			.Kernel3(32'b10111101001111001001011110100000),
			.Kernel4(32'b10111110001101101100000111100101),
			.Kernel5(32'b10111100001000110000100010011110),
			.Kernel6(32'b10111111001010101000110110101000),
			.Kernel7(32'b10111111001101011011001110011010),
			.Kernel8(32'b10111111001011011110110110100001),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*15-1:DATA_WIDHT*14]),
			.Valid_Out(CHANNEL15_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL16 (
			.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
			.Kernel0(32'b00111101100110111110101001000000),
			.Kernel1(32'b10111101100001000000000101111011),
			.Kernel2(32'b10111110100000110110011011110011),
			.Kernel3(32'b00111110100111101110010010100101),
			.Kernel4(32'b00111101001011110101001011101001),
			.Kernel5(32'b00111110110101001111101001100000),
			.Kernel6(32'b00111111001010111000110100011110),
			.Kernel7(32'b00111101110010010101000101101001),
			.Kernel8(32'b00111110101010010100100010000010),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*16-1:DATA_WIDHT*15]),
			.Valid_Out(CHANNEL16_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL17 (
			.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
			.Kernel0(32'b10111111011010000100111110011011),
			.Kernel1(32'b10111111000110101001001001100111),
			.Kernel2(32'b10111111101000011001011100101100),
			.Kernel3(32'b00111110100100111011100111101110),
			.Kernel4(32'b00111110010010011110100011000111),
			.Kernel5(32'b10111110001010101000000110111101),
			.Kernel6(32'b00111110001100001001010000011100),
			.Kernel7(32'b00111110100111011010001101010000),
			.Kernel8(32'b00111101011011000000111011110000),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*17-1:DATA_WIDHT*16]),
			.Valid_Out(CHANNEL17_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL18 (
			.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
			.Kernel0(32'b00111111010011011111000010000101),
			.Kernel1(32'b00111111010000001100110011111001),
			.Kernel2(32'b00111111010101000101101110101001),
			.Kernel3(32'b10111101100010111111001011001101),
			.Kernel4(32'b00111101010001011100110101111000),
			.Kernel5(32'b10111101000101001000010101000101),
			.Kernel6(32'b10111110111110110010001001101011),
			.Kernel7(32'b10111111000100001100100111111100),
			.Kernel8(32'b10111111000001101000111011000110),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*18-1:DATA_WIDHT*17]),
			.Valid_Out(CHANNEL18_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL19 (
			.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
			.Kernel0(32'b00111110010111000011111111111110),
			.Kernel1(32'b00111111000011010001000110000111),
			.Kernel2(32'b00111111000010100110100011001101),
			.Kernel3(32'b00111110011010110101110110101101),
			.Kernel4(32'b00111110111000101100101000011100),
			.Kernel5(32'b00111111000010110001011011101011),
			.Kernel6(32'b00111110100100001010010010011011),
			.Kernel7(32'b00111110100000111110101100100100),
			.Kernel8(32'b00111110110011000100111011111000),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*19-1:DATA_WIDHT*18]),
			.Valid_Out(CHANNEL19_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL20 (
			.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
			.Kernel0(32'b10111110100000100110011111011110),
			.Kernel1(32'b00111101111001111000100011010001),
			.Kernel2(32'b10111010011011111000001001101000),
			.Kernel3(32'b10111110101111100001110011011111),
			.Kernel4(32'b10111110101111001011001010001110),
			.Kernel5(32'b10111110111110111100110011011110),
			.Kernel6(32'b10111111000111000111110010010010),
			.Kernel7(32'b10111110000011110011011110110110),
			.Kernel8(32'b10111111001011000011000010001100),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*20-1:DATA_WIDHT*19]),
			.Valid_Out(CHANNEL20_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL21 (
			.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
			.Kernel0(32'b10111110010111000001010001001000),
			.Kernel1(32'b10111100001111101100000110000011),
			.Kernel2(32'b10111110010100111111001010110110),
			.Kernel3(32'b10111110000000011111111011011101),
			.Kernel4(32'b10111110011110011000001001001000),
			.Kernel5(32'b10111100111011000001001111001110),
			.Kernel6(32'b10111110110001011001101111100101),
			.Kernel7(32'b10111110001101110000101011110101),
			.Kernel8(32'b10111111001010100111110000111100),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*21-1:DATA_WIDHT*20]),
			.Valid_Out(CHANNEL21_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL22 (
			.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
			.Kernel0(32'b00111111001110111011001111000011),
			.Kernel1(32'b00111110111110111111011000001111),
			.Kernel2(32'b00111111000000010010010101000101),
			.Kernel3(32'b10111110011100100100111010011101),
			.Kernel4(32'b10111101110111000010001101111110),
			.Kernel5(32'b00111110100101011101101010111000),
			.Kernel6(32'b10111111011010101010001011111001),
			.Kernel7(32'b10111110100111101011000011101011),
			.Kernel8(32'b10111111001000001101000101111010),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*22-1:DATA_WIDHT*21]),
			.Valid_Out(CHANNEL22_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL23 (
			.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
			.Kernel0(32'b00111110011100001111010101011001),
			.Kernel1(32'b00111110011111000111110011110100),
			.Kernel2(32'b00111110110101011111001001101010),
			.Kernel3(32'b10111100001010000000000001110001),
			.Kernel4(32'b00111010111110001010001001010101),
			.Kernel5(32'b10111110000011010000110101010000),
			.Kernel6(32'b10111111000010001101011000111101),
			.Kernel7(32'b10111110101010001100001011110111),
			.Kernel8(32'b10111110111100001001111000101110),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*23-1:DATA_WIDHT*22]),
			.Valid_Out(CHANNEL23_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL24 (
			.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
			.Kernel0(32'b10111110101110000011110100100101),
			.Kernel1(32'b10111111001110110110000100001101),
			.Kernel2(32'b10111111010011011010101101000110),
			.Kernel3(32'b00111100010110000001001011000110),
			.Kernel4(32'b10111110100010110101111011001111),
			.Kernel5(32'b10111110111011001110111000010110),
			.Kernel6(32'b10111100110010111010111000110110),
			.Kernel7(32'b00111011010110100000010101100111),
			.Kernel8(32'b10111110100010101000101011111011),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*24-1:DATA_WIDHT*23]),
			.Valid_Out(CHANNEL24_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL25 (
			.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
			.Kernel0(32'b10111110110100101100100000100010),
			.Kernel1(32'b10111110100000110011101010011001),
			.Kernel2(32'b10111101111101101000111001010011),
			.Kernel3(32'b10111110111111001011111010111000),
			.Kernel4(32'b10111111000011111110110111011100),
			.Kernel5(32'b10111110011110011011101000011101),
			.Kernel6(32'b10111111000011011001100101111110),
			.Kernel7(32'b10111110100101101000100000101101),
			.Kernel8(32'b10111110011001011010111011100010),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*25-1:DATA_WIDHT*24]),
			.Valid_Out(CHANNEL25_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL26 (
			.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
			.Kernel0(32'b10111111000110001011001111000011),
			.Kernel1(32'b10111110110111111101010110111010),
			.Kernel2(32'b10111111011101101101110101001111),
			.Kernel3(32'b00111110001111110000110111111111),
			.Kernel4(32'b10111110011111111101110100001100),
			.Kernel5(32'b10111111001100011010110001100011),
			.Kernel6(32'b00111110110000101101100101101001),
			.Kernel7(32'b00111110001100100011001101001011),
			.Kernel8(32'b10111110011110011111010001101011),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*26-1:DATA_WIDHT*25]),
			.Valid_Out(CHANNEL26_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL27 (
			.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
			.Kernel0(32'b10111101010010101100101011001000),
			.Kernel1(32'b10111110011101100000011100010001),
			.Kernel2(32'b10111110110100100110001010010101),
			.Kernel3(32'b10111110111001101101111110001110),
			.Kernel4(32'b10111110010010010101101111001100),
			.Kernel5(32'b10111111001000110100100011011110),
			.Kernel6(32'b10111110111000010100101000100101),
			.Kernel7(32'b10111110100101100111110001011110),
			.Kernel8(32'b10111110000000010100010000001011),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*27-1:DATA_WIDHT*26]),
			.Valid_Out(CHANNEL27_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL28 (
			.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
			.Kernel0(32'b00111111000101011101111001100011),
			.Kernel1(32'b00111111001001010101101111010011),
			.Kernel2(32'b00111111001100100011001100010001),
			.Kernel3(32'b10111101110001111101010110000001),
			.Kernel4(32'b10111110111111011001111100011011),
			.Kernel5(32'b10111110101110111001001100101111),
			.Kernel6(32'b10111111001111000000110110101010),
			.Kernel7(32'b10111110111010111001010101010110),
			.Kernel8(32'b10111111000010110110001010110001),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*28-1:DATA_WIDHT*27]),
			.Valid_Out(CHANNEL28_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL29 (
			.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
			.Kernel0(32'b00111111000010001100000000000001),
			.Kernel1(32'b00111110010001101001001000101111),
			.Kernel2(32'b00111111010000110100100111110011),
			.Kernel3(32'b00111101101011101011101110010100),
			.Kernel4(32'b10111110000000110111001010100110),
			.Kernel5(32'b00111110110100110101001101010111),
			.Kernel6(32'b10111110111101010010001011000111),
			.Kernel7(32'b10111101110000001100111011101111),
			.Kernel8(32'b00111110111000010101101001010011),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*29-1:DATA_WIDHT*28]),
			.Valid_Out(CHANNEL29_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL30 (
			.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
			.Kernel0(32'b10111110111000101011110111111001),
			.Kernel1(32'b10111110001111100000000101111011),
			.Kernel2(32'b10111101011011011010110110110011),
			.Kernel3(32'b10111111000000110001100100011000),
			.Kernel4(32'b10111110011010011010111011101110),
			.Kernel5(32'b10111110100010110110111100000000),
			.Kernel6(32'b10111110010001001111101111101011),
			.Kernel7(32'b10111111000110010000000101000110),
			.Kernel8(32'b10111111001101100101011010100010),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*30-1:DATA_WIDHT*29]),
			.Valid_Out(CHANNEL30_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL31 (
			.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
			.Kernel0(32'b10111111011101010100111111001001),
			.Kernel1(32'b10111111011011011000000101100100),
			.Kernel2(32'b10111111001111010000001100101001),
			.Kernel3(32'b00111110110001101000111011001000),
			.Kernel4(32'b10111011000110010010101000000000),
			.Kernel5(32'b00111110001010111000000101011111),
			.Kernel6(32'b00111110111111100100100101110010),
			.Kernel7(32'b00111110111100100000010100100001),
			.Kernel8(32'b00111110100011001010100010110100),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*31-1:DATA_WIDHT*30]),
			.Valid_Out(CHANNEL31_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL32 (
			.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
			.Kernel0(32'b00111101010111101101011011010110),
			.Kernel1(32'b00111110010001101101110010101001),
			.Kernel2(32'b00111110111010010111011111000011),
			.Kernel3(32'b00111101111110010011010000110010),
			.Kernel4(32'b10111110100000001110001110100011),
			.Kernel5(32'b00111110000101000011111000111010),
			.Kernel6(32'b00111110011110010011010000100001),
			.Kernel7(32'b00111110100010010010110000101110),
			.Kernel8(32'b00111111000111010100001100111111),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*32-1:DATA_WIDHT*31]),
			.Valid_Out(CHANNEL32_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL33 (
			.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
			.Kernel0(32'b00111110111000000011011101110000),
			.Kernel1(32'b00111110101110010011101001000100),
			.Kernel2(32'b00111110110000111111000100110110),
			.Kernel3(32'b10111110111010011011010000010110),
			.Kernel4(32'b10111110110011000100111111001000),
			.Kernel5(32'b10111111000000111101100010110100),
			.Kernel6(32'b10111111000100001000010010101001),
			.Kernel7(32'b10111110101000010010100110101011),
			.Kernel8(32'b10111111000110001000101100111100),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*33-1:DATA_WIDHT*32]),
			.Valid_Out(CHANNEL33_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL34 (
			.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
			.Kernel0(32'b10111111000111101001010010000001),
			.Kernel1(32'b10111111000010100011100011001011),
			.Kernel2(32'b10111110111111110100100110101110),
			.Kernel3(32'b10111110001000111011000000011000),
			.Kernel4(32'b10111110100101100011101101000010),
			.Kernel5(32'b10111101110110100100111001110011),
			.Kernel6(32'b00111111001011001011101101001010),
			.Kernel7(32'b00111111000010010011010011100001),
			.Kernel8(32'b00111111000110011000110010000010),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*34-1:DATA_WIDHT*33]),
			.Valid_Out(CHANNEL34_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL35 (
			.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
			.Kernel0(32'b00111110101100111000100001010010),
			.Kernel1(32'b00111110110110110011001011001111),
			.Kernel2(32'b00111110101101000101110000010110),
			.Kernel3(32'b00111110001101010000011001110011),
			.Kernel4(32'b00111101101100100111110000000110),
			.Kernel5(32'b00111110010010111001111010101101),
			.Kernel6(32'b10111101000011111000101101001011),
			.Kernel7(32'b10111101000101001010110011101101),
			.Kernel8(32'b00111101111001101000101110110111),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*35-1:DATA_WIDHT*34]),
			.Valid_Out(CHANNEL35_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL36 (
			.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
			.Kernel0(32'b10111111000101100101100011111100),
			.Kernel1(32'b10111110111001010100010000011111),
			.Kernel2(32'b10111110011010011101110100001100),
			.Kernel3(32'b10111101110010011110101010010110),
			.Kernel4(32'b10111110000111001011010001011001),
			.Kernel5(32'b00111101010010000000111101101011),
			.Kernel6(32'b00111111001111011010100101111100),
			.Kernel7(32'b00111110101001100111001101000100),
			.Kernel8(32'b00111111000101011000111100111100),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*36-1:DATA_WIDHT*35]),
			.Valid_Out(CHANNEL36_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL37 (
			.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
			.Kernel0(32'b10111111001011000100000101011000),
			.Kernel1(32'b10111111000101110100001110110010),
			.Kernel2(32'b10111110111011000101000011100000),
			.Kernel3(32'b10111110100011000001101010111000),
			.Kernel4(32'b10111110000001000111101110000110),
			.Kernel5(32'b10111110010101001111110111100010),
			.Kernel6(32'b10111110100110010101000011000100),
			.Kernel7(32'b00111110010111101111110011110101),
			.Kernel8(32'b10111101110001101010000111100100),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*37-1:DATA_WIDHT*36]),
			.Valid_Out(CHANNEL37_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL38 (
			.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
			.Kernel0(32'b00111111011011000110110111000100),
			.Kernel1(32'b00111110100001110000010111010000),
			.Kernel2(32'b00111100101110000000001110101111),
			.Kernel3(32'b00111111010000101101111111101110),
			.Kernel4(32'b10111101001010011000001001111101),
			.Kernel5(32'b10111101000010011110010000001111),
			.Kernel6(32'b00111110111111100011011100110110),
			.Kernel7(32'b00111110010000001010000101110100),
			.Kernel8(32'b10111101101100011000011010100111),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*38-1:DATA_WIDHT*37]),
			.Valid_Out(CHANNEL38_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL39 (
			.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
			.Kernel0(32'b00111110101111101000100101101100),
			.Kernel1(32'b00111110110111110101100110100001),
			.Kernel2(32'b00111111000100101101110010111011),
			.Kernel3(32'b00111101110100111011110100110011),
			.Kernel4(32'b00111101010100100100000000011000),
			.Kernel5(32'b00111110100010011100000100100010),
			.Kernel6(32'b00111110101110001111100011110001),
			.Kernel7(32'b00111110100111100010100101010101),
			.Kernel8(32'b00111110111001011110000101100110),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*39-1:DATA_WIDHT*38]),
			.Valid_Out(CHANNEL39_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL40 (
			.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
			.Kernel0(32'b10111110000001001010110011001011),
			.Kernel1(32'b10111110001000000001001111001001),
			.Kernel2(32'b00111101101100001111011100110111),
			.Kernel3(32'b10111110010001011111111011011000),
			.Kernel4(32'b10111110000011000111101000110000),
			.Kernel5(32'b10111110101011110000011101101000),
			.Kernel6(32'b10111110111010001111011110001110),
			.Kernel7(32'b10111111000000011000100110001011),
			.Kernel8(32'b10111110111000111011000101000100),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*40-1:DATA_WIDHT*39]),
			.Valid_Out(CHANNEL40_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL41 (
			.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
			.Kernel0(32'b00111110110000000111110100100101),
			.Kernel1(32'b00111110110101001011101010101101),
			.Kernel2(32'b00111111001011101101010001001110),
			.Kernel3(32'b10111110010011000010001010001101),
			.Kernel4(32'b00111110010011001101010110101000),
			.Kernel5(32'b00111010001110111111010010001010),
			.Kernel6(32'b10111110101000100110101011110100),
			.Kernel7(32'b10111101101100010101111111101111),
			.Kernel8(32'b10111111001010001101101100101000),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*41-1:DATA_WIDHT*40]),
			.Valid_Out(CHANNEL41_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL42 (
			.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
			.Kernel0(32'b10111110011111000110001110011110),
			.Kernel1(32'b00111101110111010100000101001011),
			.Kernel2(32'b10111110111100111100011110100111),
			.Kernel3(32'b10111110001010100101110110101111),
			.Kernel4(32'b10111101001001010110011100111011),
			.Kernel5(32'b10111111001001100100000011000111),
			.Kernel6(32'b10111110101010111100100001111011),
			.Kernel7(32'b10111110101000100101000100100100),
			.Kernel8(32'b10111111000001011000000001001011),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*42-1:DATA_WIDHT*41]),
			.Valid_Out(CHANNEL42_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL43 (
			.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
			.Kernel0(32'b10111111000100110111011011011000),
			.Kernel1(32'b10111111000100000110110001100001),
			.Kernel2(32'b10111110110010100111000100100101),
			.Kernel3(32'b10111111000010111001110000010010),
			.Kernel4(32'b10111110111101001011011001101011),
			.Kernel5(32'b10111110011011010111001100011011),
			.Kernel6(32'b10111110011000010111001000100100),
			.Kernel7(32'b10111110100010000010101110101000),
			.Kernel8(32'b10111110000110100111101011110011),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*43-1:DATA_WIDHT*42]),
			.Valid_Out(CHANNEL43_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL44 (
			.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
			.Kernel0(32'b10111111000000100111101001101000),
			.Kernel1(32'b10111110100010100110011011111110),
			.Kernel2(32'b10111110110110110101111110100111),
			.Kernel3(32'b00111101111010100011001100100010),
			.Kernel4(32'b10111101110101000100000101010101),
			.Kernel5(32'b10111101111100110110111010110101),
			.Kernel6(32'b10111111000110001111001101100111),
			.Kernel7(32'b10111110100010110011010001111110),
			.Kernel8(32'b10111110110100010010101101101000),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*44-1:DATA_WIDHT*43]),
			.Valid_Out(CHANNEL44_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL45 (
			.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
			.Kernel0(32'b10111111000101110000101111000010),
			.Kernel1(32'b10111110110001100101010101110100),
			.Kernel2(32'b10111111010110100011010011011110),
			.Kernel3(32'b10111111000000000111011001011000),
			.Kernel4(32'b10111111000010111100100101011011),
			.Kernel5(32'b10111111010001011100100110110110),
			.Kernel6(32'b10111110100111111000110101011111),
			.Kernel7(32'b10111110010101100010101001100100),
			.Kernel8(32'b10111110101100001110111110110111),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*45-1:DATA_WIDHT*44]),
			.Valid_Out(CHANNEL45_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL46 (
			.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
			.Kernel0(32'b10111101100011011100100100010000),
			.Kernel1(32'b00111110010010101011111111101011),
			.Kernel2(32'b00111110101110001110011001010010),
			.Kernel3(32'b00111110100111100001010110111100),
			.Kernel4(32'b00111101101001010111110010000101),
			.Kernel5(32'b00111111001001110110001111000000),
			.Kernel6(32'b10111110100011010100010010101000),
			.Kernel7(32'b10111110011111110101101010110101),
			.Kernel8(32'b00111101101010000100100011110010),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*46-1:DATA_WIDHT*45]),
			.Valid_Out(CHANNEL46_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL47 (
			.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
			.Kernel0(32'b00111110111110111110001101110000),
			.Kernel1(32'b00111110101111000001110111010100),
			.Kernel2(32'b00111110010100101010111111101001),
			.Kernel3(32'b00111111000010100001101101101000),
			.Kernel4(32'b00111101100100110110000001111010),
			.Kernel5(32'b00111110111000001111110001111110),
			.Kernel6(32'b00111111001101101001100010110111),
			.Kernel7(32'b00111110100111000111000111101011),
			.Kernel8(32'b00111110100001010011110010000110),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*47-1:DATA_WIDHT*46]),
			.Valid_Out(CHANNEL47_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL48 (
			.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
			.Kernel0(32'b00111110111001101111110100001101),
			.Kernel1(32'b00111110100001010000110010011101),
			.Kernel2(32'b00111110110000110000100101001101),
			.Kernel3(32'b00111110110110000010010010000001),
			.Kernel4(32'b00111111000100100000011011000000),
			.Kernel5(32'b00111111010000111010000101001011),
			.Kernel6(32'b00111111011000101001010101100111),
			.Kernel7(32'b00111111001010111011111101101111),
			.Kernel8(32'b00111111001100101110000111001000),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*48-1:DATA_WIDHT*47]),
			.Valid_Out(CHANNEL48_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL49 (
			.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
			.Kernel0(32'b10111110011101101010111101100011),
			.Kernel1(32'b10111110111011101001000001110111),
			.Kernel2(32'b10111110101111111100100000110001),
			.Kernel3(32'b10111110010100110000011001001001),
			.Kernel4(32'b10111110111101111100000011000000),
			.Kernel5(32'b10111110100110011000010110001001),
			.Kernel6(32'b00111110000001010010000101101100),
			.Kernel7(32'b00111101110100011110000010101001),
			.Kernel8(32'b10111111001101000001001000101101),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*49-1:DATA_WIDHT*48]),
			.Valid_Out(CHANNEL49_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL50 (
			.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
			.Kernel0(32'b00111101100000010101010110111101),
			.Kernel1(32'b10111110100011000101110100101100),
			.Kernel2(32'b00111101100000011101100011000111),
			.Kernel3(32'b10111111000001010111010000000110),
			.Kernel4(32'b10111111000000100111100000101100),
			.Kernel5(32'b10111100010100110001001110100010),
			.Kernel6(32'b10111110111010011110101001111101),
			.Kernel7(32'b10111110110110000111111011100110),
			.Kernel8(32'b10111110100110000000110010111010),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*50-1:DATA_WIDHT*49]),
			.Valid_Out(CHANNEL50_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL51 (
			.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
			.Kernel0(32'b10111111010011011110011101101101),
			.Kernel1(32'b10111110110000000010110011001110),
			.Kernel2(32'b10111111001010100111011000011011),
			.Kernel3(32'b00111110101000100101000101001101),
			.Kernel4(32'b00111110011100100100101001010110),
			.Kernel5(32'b00111110100010001011101101000101),
			.Kernel6(32'b00111110101000001110001000010101),
			.Kernel7(32'b00111110101001100001000100010101),
			.Kernel8(32'b00111110100110001000111011010100),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*51-1:DATA_WIDHT*50]),
			.Valid_Out(CHANNEL51_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL52 (
			.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
			.Kernel0(32'b10111111000001010001101010101100),
			.Kernel1(32'b10111111000001101010001100010010),
			.Kernel2(32'b10111110100111000100010000010011),
			.Kernel3(32'b10111110000111111001000001111000),
			.Kernel4(32'b00111100100001100110010100100110),
			.Kernel5(32'b00111110000010010110010001101110),
			.Kernel6(32'b00111111000011111010111000111111),
			.Kernel7(32'b00111110111000000011000101110000),
			.Kernel8(32'b00111110111011001100100100111111),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*52-1:DATA_WIDHT*51]),
			.Valid_Out(CHANNEL52_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL53 (
			.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
			.Kernel0(32'b10111100110111011010101000010110),
			.Kernel1(32'b10111101101101110001101011101101),
			.Kernel2(32'b10111110000011110100101001110001),
			.Kernel3(32'b10111110111100111111110110011010),
			.Kernel4(32'b10111111000101000110110000011001),
			.Kernel5(32'b10111111000011001000011110100101),
			.Kernel6(32'b10111110101111000111010001111010),
			.Kernel7(32'b10111110100000011110000000101100),
			.Kernel8(32'b10111111000011101000000100001001),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*53-1:DATA_WIDHT*52]),
			.Valid_Out(CHANNEL53_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL54 (
			.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
			.Kernel0(32'b10111110100010110001111101100100),
			.Kernel1(32'b10111110110001001111101110100110),
			.Kernel2(32'b10111110110110001010110010100001),
			.Kernel3(32'b10111110110000011001011011111011),
			.Kernel4(32'b10111110010010000000010001101110),
			.Kernel5(32'b10111110100110101010111111010011),
			.Kernel6(32'b10111110110011010001111110011110),
			.Kernel7(32'b10111110110000010000000011001001),
			.Kernel8(32'b10111110100110100111011010111000),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*54-1:DATA_WIDHT*53]),
			.Valid_Out(CHANNEL54_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL55 (
			.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
			.Kernel0(32'b00111110100001110111010010001001),
			.Kernel1(32'b00111110110010011010010111000000),
			.Kernel2(32'b00111111001101001010011011100011),
			.Kernel3(32'b00111101010111110011000111001101),
			.Kernel4(32'b00111110011110111100001000110110),
			.Kernel5(32'b00111110111111100011101111110100),
			.Kernel6(32'b10111111000101001111110100000101),
			.Kernel7(32'b10111110111001110100000100000100),
			.Kernel8(32'b10111101101111101110011110011010),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*55-1:DATA_WIDHT*54]),
			.Valid_Out(CHANNEL55_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL56 (
			.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
			.Kernel0(32'b00111111010100110100100111100001),
			.Kernel1(32'b00111111010000101101001011101000),
			.Kernel2(32'b00111110010000111011110001111111),
			.Kernel3(32'b00111110111001101010111001010010),
			.Kernel4(32'b10111110100000010001100111111100),
			.Kernel5(32'b10111111000100011000010001101100),
			.Kernel6(32'b10111110100110001110010110001110),
			.Kernel7(32'b10111101000110010101010000000011),
			.Kernel8(32'b10111110101010010101000001111111),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*56-1:DATA_WIDHT*55]),
			.Valid_Out(CHANNEL56_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL57 (
			.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
			.Kernel0(32'b10111110110001011101011101000011),
			.Kernel1(32'b10111110011001001100111111100000),
			.Kernel2(32'b10111110010101011000111000000110),
			.Kernel3(32'b10111111000101110111000101010011),
			.Kernel4(32'b10111110001011111010000010110100),
			.Kernel5(32'b10111111000101101100110001111101),
			.Kernel6(32'b10111111000000100110111001001011),
			.Kernel7(32'b10111110110011010010010100010100),
			.Kernel8(32'b10111110101000111110111010010011),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*57-1:DATA_WIDHT*56]),
			.Valid_Out(CHANNEL57_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL58 (
			.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
			.Kernel0(32'b10111110100100101101111001011011),
			.Kernel1(32'b10111110001101110000110011010101),
			.Kernel2(32'b10111111010100100101000001011101),
			.Kernel3(32'b00111110111101010000110010110001),
			.Kernel4(32'b10111110010011101011101100111000),
			.Kernel5(32'b10111110001000100100011000011111),
			.Kernel6(32'b00111111000011010011101001101000),
			.Kernel7(32'b00111101001111110111100010111100),
			.Kernel8(32'b10111110101100010111110101010111),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*58-1:DATA_WIDHT*57]),
			.Valid_Out(CHANNEL58_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL59 (
			.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
			.Kernel0(32'b10111111010001000001000011001101),
			.Kernel1(32'b10111110100110010000000011000111),
			.Kernel2(32'b10111111000011100100000111011001),
			.Kernel3(32'b00111110010111000110011111100001),
			.Kernel4(32'b10111101101100010010000101001001),
			.Kernel5(32'b10111110101100010001110111101010),
			.Kernel6(32'b00111111001101110001000110110000),
			.Kernel7(32'b00111110110101011011010011101110),
			.Kernel8(32'b00111111000010111100001110000011),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*59-1:DATA_WIDHT*58]),
			.Valid_Out(CHANNEL59_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL60 (
			.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
			.Kernel0(32'b00111111010000000110110011010101),
			.Kernel1(32'b00111110100110001110100111011100),
			.Kernel2(32'b00111100111101100011011101010110),
			.Kernel3(32'b00111110111011010110101101001001),
			.Kernel4(32'b00111110000011100110010101100010),
			.Kernel5(32'b00111110100101010001100001101011),
			.Kernel6(32'b00111110111010010000111001101001),
			.Kernel7(32'b00111110110101000000011000000011),
			.Kernel8(32'b00111110100000100001011110011010),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*60-1:DATA_WIDHT*59]),
			.Valid_Out(CHANNEL60_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL61 (
			.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
			.Kernel0(32'b00111111010100101111011000100111),
			.Kernel1(32'b00111110100001101010000100000001),
			.Kernel2(32'b00111110011111000011001011110011),
			.Kernel3(32'b00111110101001011101001100110111),
			.Kernel4(32'b00111110111100010010111101001100),
			.Kernel5(32'b00111111001110100101110010000000),
			.Kernel6(32'b00111101101101110001000000101101),
			.Kernel7(32'b10111011101111001101110010111101),
			.Kernel8(32'b00111110110011011111001101001000),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*61-1:DATA_WIDHT*60]),
			.Valid_Out(CHANNEL61_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL62 (
			.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
			.Kernel0(32'b00111110100011000110110100100011),
			.Kernel1(32'b00111110101011100101101010100000),
			.Kernel2(32'b00111110011000010100100100001010),
			.Kernel3(32'b10111101101010011001111100111010),
			.Kernel4(32'b00111100110110100111010011110110),
			.Kernel5(32'b00111110001010111100110000110101),
			.Kernel6(32'b00111101000011010110010011101001),
			.Kernel7(32'b00111110101001000010110011101001),
			.Kernel8(32'b10111101101011001101110000001110),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*62-1:DATA_WIDHT*61]),
			.Valid_Out(CHANNEL62_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL63 (
			.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
			.Kernel0(32'b10111101110011101101000100001100),
			.Kernel1(32'b10111110101111010110100101101111),
			.Kernel2(32'b10111110000101100100110010100010),
			.Kernel3(32'b10111110001000010000100100101000),
			.Kernel4(32'b10111110100101111001001010101111),
			.Kernel5(32'b10111110111111110100100101100100),
			.Kernel6(32'b10111111000001111100010101000100),
			.Kernel7(32'b10111111001100001001100011110010),
			.Kernel8(32'b10111110000110110100011110111000),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*63-1:DATA_WIDHT*62]),
			.Valid_Out(CHANNEL63_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL64 (
			.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
			.Kernel0(32'b10111110110001110110001011101100),
			.Kernel1(32'b00111101011010110101011010010110),
			.Kernel2(32'b10111110100001101101010101111011),
			.Kernel3(32'b10111110110111001100101100100110),
			.Kernel4(32'b10111101101010001110001001010000),
			.Kernel5(32'b10111110101000110001100011101000),
			.Kernel6(32'b10111101011100101110110010010011),
			.Kernel7(32'b00111110000011101100101010111100),
			.Kernel8(32'b10111110011110011000000100111000),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*64-1:DATA_WIDHT*63]),
			.Valid_Out(CHANNEL64_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL65 (
			.Data_In(Data_In[DATA_WIDHT*65-1:DATA_WIDHT*64]),
			.Kernel0(32'b10111100011101111011110100101101),
			.Kernel1(32'b00111101011110111110000000000000),
			.Kernel2(32'b00111110011100011100101011111011),
			.Kernel3(32'b00111110110001001011000111100000),
			.Kernel4(32'b00111110011001000001000100100110),
			.Kernel5(32'b00111111000100001101011101011101),
			.Kernel6(32'b00111111011100011010010011101011),
			.Kernel7(32'b00111111001011000100100011100001),
			.Kernel8(32'b00111111100001111101000001000100),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*65-1:DATA_WIDHT*64]),
			.Valid_Out(CHANNEL65_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL66 (
			.Data_In(Data_In[DATA_WIDHT*66-1:DATA_WIDHT*65]),
			.Kernel0(32'b00111110101010001010010010110001),
			.Kernel1(32'b00111110100110100001110100010100),
			.Kernel2(32'b00111111001111000001001100000110),
			.Kernel3(32'b10111110101001001011010101100110),
			.Kernel4(32'b10111110001111011110101010101101),
			.Kernel5(32'b10111110010011100000110001100011),
			.Kernel6(32'b10111110111000001011110010101010),
			.Kernel7(32'b10111111000011000100001111110010),
			.Kernel8(32'b10111111001001110110111000001011),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*66-1:DATA_WIDHT*65]),
			.Valid_Out(CHANNEL66_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL67 (
			.Data_In(Data_In[DATA_WIDHT*67-1:DATA_WIDHT*66]),
			.Kernel0(32'b00111110101011100101100000111110),
			.Kernel1(32'b10111101001101110010100100001111),
			.Kernel2(32'b00111110101111100110111100111001),
			.Kernel3(32'b00111110100001010101010000111101),
			.Kernel4(32'b00111110000001010011001001110011),
			.Kernel5(32'b00111110011111101010110011101000),
			.Kernel6(32'b00111110110011101111001100001010),
			.Kernel7(32'b00111011101000111010011100111110),
			.Kernel8(32'b00111110001000000101011110010101),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*67-1:DATA_WIDHT*66]),
			.Valid_Out(CHANNEL67_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL68 (
			.Data_In(Data_In[DATA_WIDHT*68-1:DATA_WIDHT*67]),
			.Kernel0(32'b00111101110110101000000011000110),
			.Kernel1(32'b00111100110110101001011010111110),
			.Kernel2(32'b00111110011101111101010001101001),
			.Kernel3(32'b00111100111111110110100001011101),
			.Kernel4(32'b00111110001010001111011111010001),
			.Kernel5(32'b00111110100001101111111001001100),
			.Kernel6(32'b00111111000001010101000001100111),
			.Kernel7(32'b00111110111001001101100100011111),
			.Kernel8(32'b00111111000111011010011010111011),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*68-1:DATA_WIDHT*67]),
			.Valid_Out(CHANNEL68_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL69 (
			.Data_In(Data_In[DATA_WIDHT*69-1:DATA_WIDHT*68]),
			.Kernel0(32'b10111110110101000011111111111110),
			.Kernel1(32'b00111110011100100110000000000011),
			.Kernel2(32'b00111111001101001110100111111000),
			.Kernel3(32'b10111110100111001100010001000110),
			.Kernel4(32'b00111110110011101101011001100001),
			.Kernel5(32'b00111111010100000000101001110111),
			.Kernel6(32'b10111111000001110000111001111110),
			.Kernel7(32'b10111110010011011101010110001110),
			.Kernel8(32'b00111100111010001011010010011110),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*69-1:DATA_WIDHT*68]),
			.Valid_Out(CHANNEL69_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL70 (
			.Data_In(Data_In[DATA_WIDHT*70-1:DATA_WIDHT*69]),
			.Kernel0(32'b10111110110001111001100011111100),
			.Kernel1(32'b00111010100111011111110011111010),
			.Kernel2(32'b10111111000011000010010000011011),
			.Kernel3(32'b10111110100100011111010111111110),
			.Kernel4(32'b10111101100011001100011100010000),
			.Kernel5(32'b10111110110101110011000000100000),
			.Kernel6(32'b10111111000010010010101101010000),
			.Kernel7(32'b10111110000110100011100100110101),
			.Kernel8(32'b10111110011111100011100100110100),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*70-1:DATA_WIDHT*69]),
			.Valid_Out(CHANNEL70_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL71 (
			.Data_In(Data_In[DATA_WIDHT*71-1:DATA_WIDHT*70]),
			.Kernel0(32'b00111110111010000100100110000100),
			.Kernel1(32'b00111110101100010101100101000100),
			.Kernel2(32'b00111111010000100000111110101111),
			.Kernel3(32'b00111110100100111110110100111110),
			.Kernel4(32'b10111110001001000110110100001000),
			.Kernel5(32'b00111110110000110110100100110000),
			.Kernel6(32'b00111110001101110101011010011101),
			.Kernel7(32'b10111100010010110100010001110000),
			.Kernel8(32'b10111110011000010100000111101000),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*71-1:DATA_WIDHT*70]),
			.Valid_Out(CHANNEL71_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL72 (
			.Data_In(Data_In[DATA_WIDHT*72-1:DATA_WIDHT*71]),
			.Kernel0(32'b10111110100100110101001011001100),
			.Kernel1(32'b10111110101000001001110000011100),
			.Kernel2(32'b10111111000110011011001001101100),
			.Kernel3(32'b10111110000110111111010111010011),
			.Kernel4(32'b10111110101000101001000001101101),
			.Kernel5(32'b10111101110011011001101001101100),
			.Kernel6(32'b10111101111101001010111101011011),
			.Kernel7(32'b10111110101000000101100001011011),
			.Kernel8(32'b00111110010000100010100101110111),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*72-1:DATA_WIDHT*71]),
			.Valid_Out(CHANNEL72_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL73 (
			.Data_In(Data_In[DATA_WIDHT*73-1:DATA_WIDHT*72]),
			.Kernel0(32'b10111110111000101101001000111100),
			.Kernel1(32'b10111100110111110001100001101001),
			.Kernel2(32'b10111110111110101001111100100001),
			.Kernel3(32'b00111110011111110110010100011011),
			.Kernel4(32'b10111100011001000110100110000101),
			.Kernel5(32'b00111110000111100001110110111001),
			.Kernel6(32'b00111111000000111101111110011100),
			.Kernel7(32'b00111110110110001001110011110100),
			.Kernel8(32'b00111111001000110000010011001111),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*73-1:DATA_WIDHT*72]),
			.Valid_Out(CHANNEL73_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL74 (
			.Data_In(Data_In[DATA_WIDHT*74-1:DATA_WIDHT*73]),
			.Kernel0(32'b00111110000110110101111100100101),
			.Kernel1(32'b00111110110110000110001100010000),
			.Kernel2(32'b00111110101110001001001110111011),
			.Kernel3(32'b00111111000011101100001000000010),
			.Kernel4(32'b00111111001001100010100011111111),
			.Kernel5(32'b00111111001000111110001101100101),
			.Kernel6(32'b10111110110111011000101100001000),
			.Kernel7(32'b10111110100011001010001110111110),
			.Kernel8(32'b10111110101001010001010101110101),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*74-1:DATA_WIDHT*73]),
			.Valid_Out(CHANNEL74_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL75 (
			.Data_In(Data_In[DATA_WIDHT*75-1:DATA_WIDHT*74]),
			.Kernel0(32'b00111111010101111001000111011001),
			.Kernel1(32'b00111110110101000110011110010010),
			.Kernel2(32'b00111111011010100010100110011010),
			.Kernel3(32'b00111110000001101111110101111101),
			.Kernel4(32'b00111110100001000110010110100100),
			.Kernel5(32'b00111110100001010001100001010000),
			.Kernel6(32'b10111110011011001101001111011010),
			.Kernel7(32'b00111110000111111110011011101001),
			.Kernel8(32'b10111101110100110100101010001111),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*75-1:DATA_WIDHT*74]),
			.Valid_Out(CHANNEL75_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL76 (
			.Data_In(Data_In[DATA_WIDHT*76-1:DATA_WIDHT*75]),
			.Kernel0(32'b10111110001111000000010110011001),
			.Kernel1(32'b00111100101001110111000110110100),
			.Kernel2(32'b10111111000101001010110011000000),
			.Kernel3(32'b00111111000100101010100000110000),
			.Kernel4(32'b00111111000011100100011111001001),
			.Kernel5(32'b00111101100100100011001100110100),
			.Kernel6(32'b00111110111101011111101100111001),
			.Kernel7(32'b00111111010011000100011010001010),
			.Kernel8(32'b00111011010101110111000100001101),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*76-1:DATA_WIDHT*75]),
			.Valid_Out(CHANNEL76_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL77 (
			.Data_In(Data_In[DATA_WIDHT*77-1:DATA_WIDHT*76]),
			.Kernel0(32'b10111111010011101111000101001110),
			.Kernel1(32'b10111111001110100111001110100010),
			.Kernel2(32'b10111110111101010101100001000100),
			.Kernel3(32'b10111110110100101101000011101011),
			.Kernel4(32'b10111111001111010010101100100011),
			.Kernel5(32'b10111111000011110111101101101111),
			.Kernel6(32'b10111110000000110111010010110000),
			.Kernel7(32'b10111110100100010001111111101100),
			.Kernel8(32'b10111111010100111110100010010100),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*77-1:DATA_WIDHT*76]),
			.Valid_Out(CHANNEL77_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL78 (
			.Data_In(Data_In[DATA_WIDHT*78-1:DATA_WIDHT*77]),
			.Kernel0(32'b00111111000101100100000010010111),
			.Kernel1(32'b00111101100000110110010100010110),
			.Kernel2(32'b00111111000011001000101001010111),
			.Kernel3(32'b00111111000110001011011000101100),
			.Kernel4(32'b00111111000010111011110111011111),
			.Kernel5(32'b00111110111100011100111011111011),
			.Kernel6(32'b00111111000011010100000111010001),
			.Kernel7(32'b00111110011000011010100101010101),
			.Kernel8(32'b00111111000010101111111111101010),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*78-1:DATA_WIDHT*77]),
			.Valid_Out(CHANNEL78_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL79 (
			.Data_In(Data_In[DATA_WIDHT*79-1:DATA_WIDHT*78]),
			.Kernel0(32'b10111110111010110001001010110110),
			.Kernel1(32'b10111110101011111010110010110001),
			.Kernel2(32'b10111111001010000101001111000011),
			.Kernel3(32'b10111111000101011100101111111000),
			.Kernel4(32'b10111111000000001110000110110110),
			.Kernel5(32'b10111110100001101111001010000101),
			.Kernel6(32'b00111110101111001000001111111110),
			.Kernel7(32'b00111110000101011011010011011010),
			.Kernel8(32'b00111111000001000000100110100011),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*79-1:DATA_WIDHT*78]),
			.Valid_Out(CHANNEL79_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL80 (
			.Data_In(Data_In[DATA_WIDHT*80-1:DATA_WIDHT*79]),
			.Kernel0(32'b10111110110000010101011001110111),
			.Kernel1(32'b10111101110111001011111001100011),
			.Kernel2(32'b10111110011111100001000110010110),
			.Kernel3(32'b10111110110110110110001100011100),
			.Kernel4(32'b10111110010011101100001011111011),
			.Kernel5(32'b10111110101011111001001010101101),
			.Kernel6(32'b10111110010000110101100001000001),
			.Kernel7(32'b10111110100001111001100011011111),
			.Kernel8(32'b10111110111001011011000010000111),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*80-1:DATA_WIDHT*79]),
			.Valid_Out(CHANNEL80_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL81 (
			.Data_In(Data_In[DATA_WIDHT*81-1:DATA_WIDHT*80]),
			.Kernel0(32'b00111110000110111100110000101111),
			.Kernel1(32'b00111110110111110001110001110010),
			.Kernel2(32'b00111111001010001100000101000111),
			.Kernel3(32'b00111111000101010111100011101101),
			.Kernel4(32'b00111111000011110110111001110001),
			.Kernel5(32'b00111111001111111000110000001101),
			.Kernel6(32'b10111110101110010001111001100101),
			.Kernel7(32'b10111110100110100101100110110000),
			.Kernel8(32'b10111110011011110100010100100010),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*81-1:DATA_WIDHT*80]),
			.Valid_Out(CHANNEL81_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL82 (
			.Data_In(Data_In[DATA_WIDHT*82-1:DATA_WIDHT*81]),
			.Kernel0(32'b00111101111011101011100110011100),
			.Kernel1(32'b00111110010010001100110010001100),
			.Kernel2(32'b00111110100100101011001100101011),
			.Kernel3(32'b00111101101001101100011110100101),
			.Kernel4(32'b00111110101000011110110110111011),
			.Kernel5(32'b00111110100111111100010000111101),
			.Kernel6(32'b00111111001010000000100111000011),
			.Kernel7(32'b00111110111111110110010000000100),
			.Kernel8(32'b00111110110000111111000110110110),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*82-1:DATA_WIDHT*81]),
			.Valid_Out(CHANNEL82_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL83 (
			.Data_In(Data_In[DATA_WIDHT*83-1:DATA_WIDHT*82]),
			.Kernel0(32'b00111110000110011111001111001001),
			.Kernel1(32'b00111101100001010101111100101101),
			.Kernel2(32'b00111110001011111011000101001100),
			.Kernel3(32'b00111110101101101001001110111101),
			.Kernel4(32'b00111110101001011110010110101011),
			.Kernel5(32'b00111110000110110111011101001011),
			.Kernel6(32'b00111110110111101111101110001001),
			.Kernel7(32'b00111110110010111000100011001000),
			.Kernel8(32'b00111111000101111010001011001010),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*83-1:DATA_WIDHT*82]),
			.Valid_Out(CHANNEL83_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL84 (
			.Data_In(Data_In[DATA_WIDHT*84-1:DATA_WIDHT*83]),
			.Kernel0(32'b00111110100101001000001001101000),
			.Kernel1(32'b00111101101101000010101101000011),
			.Kernel2(32'b00111110010011011010100110110000),
			.Kernel3(32'b00111110011000010001110010000110),
			.Kernel4(32'b00111110001111110100111101100000),
			.Kernel5(32'b00111110100111111110100001100011),
			.Kernel6(32'b00111110101011100110101100111001),
			.Kernel7(32'b00111110100000010001010110111000),
			.Kernel8(32'b00111110011101101011111101100001),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*84-1:DATA_WIDHT*83]),
			.Valid_Out(CHANNEL84_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL85 (
			.Data_In(Data_In[DATA_WIDHT*85-1:DATA_WIDHT*84]),
			.Kernel0(32'b10111110101110110100101010100101),
			.Kernel1(32'b10111110111111100111000100010101),
			.Kernel2(32'b10111111000111010010001001110000),
			.Kernel3(32'b10111110111110010101111011000101),
			.Kernel4(32'b00111110000111001011100101111111),
			.Kernel5(32'b00111101111010101100011010110101),
			.Kernel6(32'b00111110101101010010100000000001),
			.Kernel7(32'b00111110110001010101000010110010),
			.Kernel8(32'b00111110010100000111111000110001),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*85-1:DATA_WIDHT*84]),
			.Valid_Out(CHANNEL85_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL86 (
			.Data_In(Data_In[DATA_WIDHT*86-1:DATA_WIDHT*85]),
			.Kernel0(32'b00111110101000100110111001100011),
			.Kernel1(32'b00111110101001100010010101111000),
			.Kernel2(32'b00111110011010010101010000001011),
			.Kernel3(32'b00111101111111010110100110010010),
			.Kernel4(32'b00111111000000010001010000001010),
			.Kernel5(32'b10111101000000011101100111000111),
			.Kernel6(32'b00111110111100100110011000000111),
			.Kernel7(32'b00111110110001100001011100100011),
			.Kernel8(32'b10111101001101010010001001010010),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*86-1:DATA_WIDHT*85]),
			.Valid_Out(CHANNEL86_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL87 (
			.Data_In(Data_In[DATA_WIDHT*87-1:DATA_WIDHT*86]),
			.Kernel0(32'b10111111001001100001000110100010),
			.Kernel1(32'b10111111001001001111001011001111),
			.Kernel2(32'b10111110101110011100100001111011),
			.Kernel3(32'b10111111000001111011000110110100),
			.Kernel4(32'b00111101111010001001101101010010),
			.Kernel5(32'b10111101111000010111101010010001),
			.Kernel6(32'b00111110100111110011110001011011),
			.Kernel7(32'b00111110111110110100011100110001),
			.Kernel8(32'b00111111001010010101111101111101),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*87-1:DATA_WIDHT*86]),
			.Valid_Out(CHANNEL87_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL88 (
			.Data_In(Data_In[DATA_WIDHT*88-1:DATA_WIDHT*87]),
			.Kernel0(32'b10111110101111001110011110001010),
			.Kernel1(32'b10111110110000110111100001110101),
			.Kernel2(32'b00111110001010101000100010111001),
			.Kernel3(32'b10111111000100110000101110011000),
			.Kernel4(32'b10111110111111011001110101100101),
			.Kernel5(32'b10111101010011001011011010101010),
			.Kernel6(32'b10111111000111100101100110011101),
			.Kernel7(32'b10111111001100000111110111010100),
			.Kernel8(32'b10111111000100111110011110010100),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*88-1:DATA_WIDHT*87]),
			.Valid_Out(CHANNEL88_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL89 (
			.Data_In(Data_In[DATA_WIDHT*89-1:DATA_WIDHT*88]),
			.Kernel0(32'b00111110101100010110010110100011),
			.Kernel1(32'b00111111000010010110100100101101),
			.Kernel2(32'b00111110110000010000111000010011),
			.Kernel3(32'b00111110111111010011110001100111),
			.Kernel4(32'b00111110111001001011010110110011),
			.Kernel5(32'b00111110111111110000001100110100),
			.Kernel6(32'b00111111000011100110000000001100),
			.Kernel7(32'b00111110110110011011000011011111),
			.Kernel8(32'b00111111001000000010001001000111),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*89-1:DATA_WIDHT*88]),
			.Valid_Out(CHANNEL89_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL90 (
			.Data_In(Data_In[DATA_WIDHT*90-1:DATA_WIDHT*89]),
			.Kernel0(32'b00111110100000000110100010110110),
			.Kernel1(32'b00111110110011110101000000010000),
			.Kernel2(32'b00111110101010101001011001111101),
			.Kernel3(32'b00111110100001011110101001110100),
			.Kernel4(32'b00111101110011001010111110101101),
			.Kernel5(32'b00111110111000000100111001001110),
			.Kernel6(32'b00111110101001001001001111101111),
			.Kernel7(32'b00111110001000011101111100001001),
			.Kernel8(32'b00111110001101110100001010001000),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*90-1:DATA_WIDHT*89]),
			.Valid_Out(CHANNEL90_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL91 (
			.Data_In(Data_In[DATA_WIDHT*91-1:DATA_WIDHT*90]),
			.Kernel0(32'b10111111000111100111100010110001),
			.Kernel1(32'b10111110000100110100110010010100),
			.Kernel2(32'b10111111000110100000101101111111),
			.Kernel3(32'b10111110101111110011011110110010),
			.Kernel4(32'b10111101101101011000000010001110),
			.Kernel5(32'b00111110000010100110010110000000),
			.Kernel6(32'b10111101101110001111000011001100),
			.Kernel7(32'b10111110011010010001111101001100),
			.Kernel8(32'b10111100111010000001101100101011),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*91-1:DATA_WIDHT*90]),
			.Valid_Out(CHANNEL91_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL92 (
			.Data_In(Data_In[DATA_WIDHT*92-1:DATA_WIDHT*91]),
			.Kernel0(32'b10111110000110111011001001011000),
			.Kernel1(32'b10111101111001001010110010100010),
			.Kernel2(32'b10111101110001101011110010000111),
			.Kernel3(32'b10111110111010111001001001110110),
			.Kernel4(32'b10111110110001111101101010011001),
			.Kernel5(32'b10111101101010110100110110110010),
			.Kernel6(32'b10111111000001011101000100010101),
			.Kernel7(32'b10111110111010101001100100000110),
			.Kernel8(32'b10111111001100010001100111111110),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*92-1:DATA_WIDHT*91]),
			.Valid_Out(CHANNEL92_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL93 (
			.Data_In(Data_In[DATA_WIDHT*93-1:DATA_WIDHT*92]),
			.Kernel0(32'b10111011100101100100101000111011),
			.Kernel1(32'b10111110100111001011000001011010),
			.Kernel2(32'b10111110110001011100111101100100),
			.Kernel3(32'b10111111001000101111011010110110),
			.Kernel4(32'b10111110111000100101011000100111),
			.Kernel5(32'b10111110101011101110000110100010),
			.Kernel6(32'b00111110101100001011001110110100),
			.Kernel7(32'b00111111001011111101111010000000),
			.Kernel8(32'b00111111001100101000000100101001),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*93-1:DATA_WIDHT*92]),
			.Valid_Out(CHANNEL93_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL94 (
			.Data_In(Data_In[DATA_WIDHT*94-1:DATA_WIDHT*93]),
			.Kernel0(32'b10111111001001011000100101000010),
			.Kernel1(32'b10111110110110000000111000010011),
			.Kernel2(32'b10111110111010010000000111011010),
			.Kernel3(32'b10111110001110010111101111011001),
			.Kernel4(32'b00111100111011111111001101100000),
			.Kernel5(32'b10111101011011010110111011111001),
			.Kernel6(32'b10111110100101010101100011001100),
			.Kernel7(32'b00111110000011110010001111010111),
			.Kernel8(32'b00111101100110000111000011101001),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*94-1:DATA_WIDHT*93]),
			.Valid_Out(CHANNEL94_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL95 (
			.Data_In(Data_In[DATA_WIDHT*95-1:DATA_WIDHT*94]),
			.Kernel0(32'b00111110100000000100000100111100),
			.Kernel1(32'b00111110111000000111101001100101),
			.Kernel2(32'b00111110111000101100110011111010),
			.Kernel3(32'b00111111010110110010001011100101),
			.Kernel4(32'b00111110100110100100100000110111),
			.Kernel5(32'b00111111010100010011100000001101),
			.Kernel6(32'b00111110111110111010111100101100),
			.Kernel7(32'b00111111000000011111101000000111),
			.Kernel8(32'b00111110011010001001111010100110),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*95-1:DATA_WIDHT*94]),
			.Valid_Out(CHANNEL95_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL96 (
			.Data_In(Data_In[DATA_WIDHT*96-1:DATA_WIDHT*95]),
			.Kernel0(32'b10111110100010010100000100101000),
			.Kernel1(32'b00111110001101000101110000101101),
			.Kernel2(32'b10111110101100111111011100100000),
			.Kernel3(32'b10111111010110111011000101011111),
			.Kernel4(32'b10111111001001101011010000100011),
			.Kernel5(32'b10111110110010001011110011101000),
			.Kernel6(32'b10111110110011101011100110001111),
			.Kernel7(32'b10111110101010100110111101011100),
			.Kernel8(32'b10111110111111000110010110000011),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*96-1:DATA_WIDHT*95]),
			.Valid_Out(CHANNEL96_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL97 (
			.Data_In(Data_In[DATA_WIDHT*97-1:DATA_WIDHT*96]),
			.Kernel0(32'b10111111000111111011001100001110),
			.Kernel1(32'b10111111000010000100110000010010),
			.Kernel2(32'b00111101011110000110111001001010),
			.Kernel3(32'b10111110101111101001000001101100),
			.Kernel4(32'b10111101100000100110010010011101),
			.Kernel5(32'b00111110010111100110110100100100),
			.Kernel6(32'b10111111000100000011000101000101),
			.Kernel7(32'b10111110100001001010011011011101),
			.Kernel8(32'b00111110001010010110100001001101),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*97-1:DATA_WIDHT*96]),
			.Valid_Out(CHANNEL97_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL98 (
			.Data_In(Data_In[DATA_WIDHT*98-1:DATA_WIDHT*97]),
			.Kernel0(32'b10111110111101101100101000110111),
			.Kernel1(32'b00111100011000010011110110110110),
			.Kernel2(32'b10111110100001010110001010001000),
			.Kernel3(32'b10111110111011100110010100111010),
			.Kernel4(32'b10111111000100110011101010001111),
			.Kernel5(32'b10111110111000110001010011010101),
			.Kernel6(32'b10111110110100011011001011101111),
			.Kernel7(32'b10111110111110101010011000111001),
			.Kernel8(32'b10111110100110010001001111001010),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*98-1:DATA_WIDHT*97]),
			.Valid_Out(CHANNEL98_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL99 (
			.Data_In(Data_In[DATA_WIDHT*99-1:DATA_WIDHT*98]),
			.Kernel0(32'b10111111011001000100011110101100),
			.Kernel1(32'b10111111001111001011011010111110),
			.Kernel2(32'b10111111011001110100011000010100),
			.Kernel3(32'b10111001011100111010101011101010),
			.Kernel4(32'b10111110000001011000010010111000),
			.Kernel5(32'b10111111000101010010000000101011),
			.Kernel6(32'b10111100101111110001101000111110),
			.Kernel7(32'b00111110000101110000111001101100),
			.Kernel8(32'b10111110000000001000101111011000),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*99-1:DATA_WIDHT*98]),
			.Valid_Out(CHANNEL99_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL100 (
			.Data_In(Data_In[DATA_WIDHT*100-1:DATA_WIDHT*99]),
			.Kernel0(32'b00111110010011011111000100110000),
			.Kernel1(32'b00111110000101101101111001110000),
			.Kernel2(32'b00111111000101100111100100110110),
			.Kernel3(32'b00111111000111011100111001100011),
			.Kernel4(32'b00111110111011111110001111100001),
			.Kernel5(32'b00111110000111111010101011000001),
			.Kernel6(32'b00111101111000100100000100110111),
			.Kernel7(32'b10111101010101110000010010011010),
			.Kernel8(32'b10111110000010000101101010010110),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*100-1:DATA_WIDHT*99]),
			.Valid_Out(CHANNEL100_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL101 (
			.Data_In(Data_In[DATA_WIDHT*101-1:DATA_WIDHT*100]),
			.Kernel0(32'b10111110101011111001011001001001),
			.Kernel1(32'b10111110100010111000111010011111),
			.Kernel2(32'b10111110101111101010010100111101),
			.Kernel3(32'b10111110010111101110101010111100),
			.Kernel4(32'b10111101110010101000101111110011),
			.Kernel5(32'b10111110110111010000010000000111),
			.Kernel6(32'b10111110111110000010111010001010),
			.Kernel7(32'b10111100101101101000101101101101),
			.Kernel8(32'b10111110110000101000001110100100),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*101-1:DATA_WIDHT*100]),
			.Valid_Out(CHANNEL101_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL102 (
			.Data_In(Data_In[DATA_WIDHT*102-1:DATA_WIDHT*101]),
			.Kernel0(32'b00111111001100100001000110100101),
			.Kernel1(32'b00111111001010010110100000001011),
			.Kernel2(32'b00111110011011111010100101001100),
			.Kernel3(32'b00111111000010110011010101001101),
			.Kernel4(32'b00111110101100000101001000000010),
			.Kernel5(32'b00111110110110000110100110110111),
			.Kernel6(32'b00111100100011100101111111101110),
			.Kernel7(32'b00111110111010111010010101100000),
			.Kernel8(32'b00111110010111111101100111010110),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*102-1:DATA_WIDHT*101]),
			.Valid_Out(CHANNEL102_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL103 (
			.Data_In(Data_In[DATA_WIDHT*103-1:DATA_WIDHT*102]),
			.Kernel0(32'b00111111000011001011000110001010),
			.Kernel1(32'b00111110110010001100100110110110),
			.Kernel2(32'b00111110100001111000100100000111),
			.Kernel3(32'b00111110101010001011110001111111),
			.Kernel4(32'b00111110000000100010010111101111),
			.Kernel5(32'b10111110011011101000000110111111),
			.Kernel6(32'b10111111000100000101101011100011),
			.Kernel7(32'b10111110110011011100011001101011),
			.Kernel8(32'b10111111000100010001010111110100),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*103-1:DATA_WIDHT*102]),
			.Valid_Out(CHANNEL103_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL104 (
			.Data_In(Data_In[DATA_WIDHT*104-1:DATA_WIDHT*103]),
			.Kernel0(32'b00111100001000101011000101110110),
			.Kernel1(32'b10111101110110101000100001010010),
			.Kernel2(32'b00111111000010111010110111111100),
			.Kernel3(32'b00111110100001100101110011100111),
			.Kernel4(32'b00111110101011000010011101111110),
			.Kernel5(32'b00111110110001111000011111100011),
			.Kernel6(32'b00111110001100001000011001000110),
			.Kernel7(32'b10111101011000001111000110111110),
			.Kernel8(32'b00111110001101101111100100011011),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*104-1:DATA_WIDHT*103]),
			.Valid_Out(CHANNEL104_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL105 (
			.Data_In(Data_In[DATA_WIDHT*105-1:DATA_WIDHT*104]),
			.Kernel0(32'b10111111000110011101110011100111),
			.Kernel1(32'b10111110111101101101010100100010),
			.Kernel2(32'b10111110110011100011001011101101),
			.Kernel3(32'b10111110101110001011101101001101),
			.Kernel4(32'b10111110110001101101001111111001),
			.Kernel5(32'b10111111001111011010010000011010),
			.Kernel6(32'b00111110100100101110111001111110),
			.Kernel7(32'b00111110000001110011011101001100),
			.Kernel8(32'b00111110110001000100110100100010),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*105-1:DATA_WIDHT*104]),
			.Valid_Out(CHANNEL105_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL106 (
			.Data_In(Data_In[DATA_WIDHT*106-1:DATA_WIDHT*105]),
			.Kernel0(32'b10111110010110100110001111100001),
			.Kernel1(32'b10111110011100000101110100011100),
			.Kernel2(32'b10111110110010000011001110011100),
			.Kernel3(32'b10111110111100110101110011001001),
			.Kernel4(32'b10111110111011111100101011110110),
			.Kernel5(32'b10111110101111110110000111010111),
			.Kernel6(32'b00111101110110111101001001010001),
			.Kernel7(32'b10111101101010111010000101000111),
			.Kernel8(32'b10111110011010110110111101001100),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*106-1:DATA_WIDHT*105]),
			.Valid_Out(CHANNEL106_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL107 (
			.Data_In(Data_In[DATA_WIDHT*107-1:DATA_WIDHT*106]),
			.Kernel0(32'b10111110010100001010001001110111),
			.Kernel1(32'b00111110101111001011110001011001),
			.Kernel2(32'b00111110110000111100011010010110),
			.Kernel3(32'b10111111000001000110010001111100),
			.Kernel4(32'b10111110111011010101011111011100),
			.Kernel5(32'b10111100011100111100111000000111),
			.Kernel6(32'b10111110011101101000011011111100),
			.Kernel7(32'b10111111000011001010101110000001),
			.Kernel8(32'b10111111001000010000000000000110),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*107-1:DATA_WIDHT*106]),
			.Valid_Out(CHANNEL107_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL108 (
			.Data_In(Data_In[DATA_WIDHT*108-1:DATA_WIDHT*107]),
			.Kernel0(32'b10111110010000111000010101111110),
			.Kernel1(32'b10111101101010101000100100010111),
			.Kernel2(32'b10111110110010101000011001001111),
			.Kernel3(32'b10111111001011101011100001111111),
			.Kernel4(32'b10111110101000011000111110111011),
			.Kernel5(32'b10111110111011001101011010110101),
			.Kernel6(32'b10111110111001000011000010011111),
			.Kernel7(32'b10111110011100100000000110110101),
			.Kernel8(32'b10111110010001101111001000101110),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*108-1:DATA_WIDHT*107]),
			.Valid_Out(CHANNEL108_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL109 (
			.Data_In(Data_In[DATA_WIDHT*109-1:DATA_WIDHT*108]),
			.Kernel0(32'b10111110110101101111111110011111),
			.Kernel1(32'b10111101111101011010010100011111),
			.Kernel2(32'b10111111010000011111000000000111),
			.Kernel3(32'b00111110000101101010111000010110),
			.Kernel4(32'b10111110001000100010101101011010),
			.Kernel5(32'b10111110110100110101101010101111),
			.Kernel6(32'b00111111010001010001101100111101),
			.Kernel7(32'b00111110101100010001000001011011),
			.Kernel8(32'b00111110101100111000110101111011),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*109-1:DATA_WIDHT*108]),
			.Valid_Out(CHANNEL109_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL110 (
			.Data_In(Data_In[DATA_WIDHT*110-1:DATA_WIDHT*109]),
			.Kernel0(32'b00111111001001100111100001010011),
			.Kernel1(32'b00111101101010111000110001110011),
			.Kernel2(32'b00111110000111000000110111010011),
			.Kernel3(32'b00111110110101100001010001001000),
			.Kernel4(32'b00111111001001000001100111100001),
			.Kernel5(32'b00111111000111110101010000011010),
			.Kernel6(32'b00111011111110011011100100101010),
			.Kernel7(32'b00111110001000101010110001101011),
			.Kernel8(32'b00111101011011011010010100101101),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*110-1:DATA_WIDHT*109]),
			.Valid_Out(CHANNEL110_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL111 (
			.Data_In(Data_In[DATA_WIDHT*111-1:DATA_WIDHT*110]),
			.Kernel0(32'b00111111001111011001011010101100),
			.Kernel1(32'b00111110110111001110101000010011),
			.Kernel2(32'b00111110010100111100000110111011),
			.Kernel3(32'b00111110011011010010000000000100),
			.Kernel4(32'b10111110010000101000011010111000),
			.Kernel5(32'b10111110111000001010100011011100),
			.Kernel6(32'b10111110100000000001000110101100),
			.Kernel7(32'b10111110101001010110111110111100),
			.Kernel8(32'b10111110101010101101011101010101),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*111-1:DATA_WIDHT*110]),
			.Valid_Out(CHANNEL111_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL112 (
			.Data_In(Data_In[DATA_WIDHT*112-1:DATA_WIDHT*111]),
			.Kernel0(32'b00111111010100110110001011110111),
			.Kernel1(32'b00111110100000011011111101111011),
			.Kernel2(32'b00111111000011011101101100001110),
			.Kernel3(32'b00111100111011010000101000100101),
			.Kernel4(32'b10111110001110010101100101000001),
			.Kernel5(32'b00111100101000101101001011110001),
			.Kernel6(32'b10111110110010000111110110010111),
			.Kernel7(32'b10111101111000101100110010011111),
			.Kernel8(32'b10111110100000110001010110101111),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*112-1:DATA_WIDHT*111]),
			.Valid_Out(CHANNEL112_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL113 (
			.Data_In(Data_In[DATA_WIDHT*113-1:DATA_WIDHT*112]),
			.Kernel0(32'b00111110010001001010010001001001),
			.Kernel1(32'b00111110100000111010100111010000),
			.Kernel2(32'b00111110101100110111100111010011),
			.Kernel3(32'b10111111000011000000010001011000),
			.Kernel4(32'b10111110100111011000110011000011),
			.Kernel5(32'b10111101111011110101010101111100),
			.Kernel6(32'b10111110111001000011001001101111),
			.Kernel7(32'b10111110110010010100011101111011),
			.Kernel8(32'b00111101100111110001010001001101),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*113-1:DATA_WIDHT*112]),
			.Valid_Out(CHANNEL113_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL114 (
			.Data_In(Data_In[DATA_WIDHT*114-1:DATA_WIDHT*113]),
			.Kernel0(32'b00111101101000110010101111011111),
			.Kernel1(32'b00111100111000111011100111010111),
			.Kernel2(32'b10111110100111011001110101001010),
			.Kernel3(32'b00111111000101101111110010110001),
			.Kernel4(32'b00111111000111001011100010101011),
			.Kernel5(32'b00111111001100000000011100000010),
			.Kernel6(32'b10111110001100110000100011001110),
			.Kernel7(32'b10111110000110000000100010011000),
			.Kernel8(32'b10111110010001001100001011011000),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*114-1:DATA_WIDHT*113]),
			.Valid_Out(CHANNEL114_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL115 (
			.Data_In(Data_In[DATA_WIDHT*115-1:DATA_WIDHT*114]),
			.Kernel0(32'b00111111010100011000010001100001),
			.Kernel1(32'b00111110011001011110110100000001),
			.Kernel2(32'b00111111001000100110001100001111),
			.Kernel3(32'b00111101110100010010011000011100),
			.Kernel4(32'b00111101101001111111100110100101),
			.Kernel5(32'b00111110000000010101110000011100),
			.Kernel6(32'b10111110110000100100100101001101),
			.Kernel7(32'b10111110001001100001010111001000),
			.Kernel8(32'b10111110011111101010010000000010),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*115-1:DATA_WIDHT*114]),
			.Valid_Out(CHANNEL115_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL116 (
			.Data_In(Data_In[DATA_WIDHT*116-1:DATA_WIDHT*115]),
			.Kernel0(32'b00111110101111001100101111010110),
			.Kernel1(32'b00111110011101010101101100101100),
			.Kernel2(32'b00111110000011110111111000101001),
			.Kernel3(32'b00111110110000001100111011000111),
			.Kernel4(32'b00111110111101001101010101011011),
			.Kernel5(32'b00111111000101001000101010101110),
			.Kernel6(32'b00111110110101101101011011110010),
			.Kernel7(32'b00111110111111111101110010000110),
			.Kernel8(32'b00111111000011010100010100010101),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*116-1:DATA_WIDHT*115]),
			.Valid_Out(CHANNEL116_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL117 (
			.Data_In(Data_In[DATA_WIDHT*117-1:DATA_WIDHT*116]),
			.Kernel0(32'b00111110111010101100100001001100),
			.Kernel1(32'b00111111000010010011100111010010),
			.Kernel2(32'b00111111000101101011000011010010),
			.Kernel3(32'b00111111010001001001010100110111),
			.Kernel4(32'b00111111000000011001101110011111),
			.Kernel5(32'b00111111000110111011010011000011),
			.Kernel6(32'b10111110111011100010101110100011),
			.Kernel7(32'b10111110101000111010001101111001),
			.Kernel8(32'b10111110101110100110000011100110),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*117-1:DATA_WIDHT*116]),
			.Valid_Out(CHANNEL117_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL118 (
			.Data_In(Data_In[DATA_WIDHT*118-1:DATA_WIDHT*117]),
			.Kernel0(32'b10111110111101000100010011100011),
			.Kernel1(32'b10111110001101111000111000000101),
			.Kernel2(32'b00111100101010111011000000010111),
			.Kernel3(32'b10111111000001100101110100010011),
			.Kernel4(32'b10111110011100101111011101011110),
			.Kernel5(32'b00111110000001011111100100011010),
			.Kernel6(32'b10111111001001000110100101000101),
			.Kernel7(32'b00111110101000010110001101010111),
			.Kernel8(32'b00111111001011010100110101010000),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*118-1:DATA_WIDHT*117]),
			.Valid_Out(CHANNEL118_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL119 (
			.Data_In(Data_In[DATA_WIDHT*119-1:DATA_WIDHT*118]),
			.Kernel0(32'b10111110110110010111100011010010),
			.Kernel1(32'b10111101100100111001001111001111),
			.Kernel2(32'b10111111001000011011000110000010),
			.Kernel3(32'b10111110000101100110010101100010),
			.Kernel4(32'b00111101101001000110110111100000),
			.Kernel5(32'b00111110011100001000111100101110),
			.Kernel6(32'b00111111000011011110010011100110),
			.Kernel7(32'b00111110111011100011100111110110),
			.Kernel8(32'b00111111001101010111011111101000),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*119-1:DATA_WIDHT*118]),
			.Valid_Out(CHANNEL119_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL120 (
			.Data_In(Data_In[DATA_WIDHT*120-1:DATA_WIDHT*119]),
			.Kernel0(32'b00111101110101101011100101110001),
			.Kernel1(32'b00111110010101101101111100000000),
			.Kernel2(32'b10111101111001011000001001011101),
			.Kernel3(32'b00111101101010100000101101100110),
			.Kernel4(32'b00111110101010100001100110010011),
			.Kernel5(32'b00111101110101110110101100010010),
			.Kernel6(32'b00111111000011010000101100101011),
			.Kernel7(32'b00111111001010100000101010100000),
			.Kernel8(32'b00111111001001000011100101101001),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*120-1:DATA_WIDHT*119]),
			.Valid_Out(CHANNEL120_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL121 (
			.Data_In(Data_In[DATA_WIDHT*121-1:DATA_WIDHT*120]),
			.Kernel0(32'b00111011101001100101100011010001),
			.Kernel1(32'b00111110010100010100100010111100),
			.Kernel2(32'b00111110100100010111111011110010),
			.Kernel3(32'b00111111000111101101100010100110),
			.Kernel4(32'b00111111000101111010011101001111),
			.Kernel5(32'b00111111010011100001010101100111),
			.Kernel6(32'b00111111000010000111011000101011),
			.Kernel7(32'b00111111011000111111000110000110),
			.Kernel8(32'b00111111011100000101011101111010),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*121-1:DATA_WIDHT*120]),
			.Valid_Out(CHANNEL121_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL122 (
			.Data_In(Data_In[DATA_WIDHT*122-1:DATA_WIDHT*121]),
			.Kernel0(32'b10111101110110000010010010010001),
			.Kernel1(32'b00111110001111010101011011001100),
			.Kernel2(32'b10111101001111001111010001011001),
			.Kernel3(32'b00111110100001110001001111111110),
			.Kernel4(32'b00111110110010110010111010000100),
			.Kernel5(32'b00111110010101011001011011110111),
			.Kernel6(32'b00111111001011011111111001101100),
			.Kernel7(32'b00111111000110010011110101111111),
			.Kernel8(32'b00111111000110000000100101100001),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*122-1:DATA_WIDHT*121]),
			.Valid_Out(CHANNEL122_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL123 (
			.Data_In(Data_In[DATA_WIDHT*123-1:DATA_WIDHT*122]),
			.Kernel0(32'b00111101100010001010111010001011),
			.Kernel1(32'b10111111000010010010010000101001),
			.Kernel2(32'b10111110100101101110011110011111),
			.Kernel3(32'b10111101011001111101000100010111),
			.Kernel4(32'b10111111000111000111011100110100),
			.Kernel5(32'b10111110100010100000110011010100),
			.Kernel6(32'b10111110100010000001100111110010),
			.Kernel7(32'b10111111001111101110110001110011),
			.Kernel8(32'b10111110111001101011010101001010),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*123-1:DATA_WIDHT*122]),
			.Valid_Out(CHANNEL123_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL124 (
			.Data_In(Data_In[DATA_WIDHT*124-1:DATA_WIDHT*123]),
			.Kernel0(32'b10111111010001100111111000001100),
			.Kernel1(32'b10111111001000000000101110001100),
			.Kernel2(32'b10111110101100000111001101110100),
			.Kernel3(32'b10111110100011010101111100100001),
			.Kernel4(32'b10111101001111010111100111111101),
			.Kernel5(32'b00111110011101101001101111000111),
			.Kernel6(32'b00111110111011001000010010101000),
			.Kernel7(32'b00111111001010101110100100111000),
			.Kernel8(32'b00111111000111101110010100010101),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*124-1:DATA_WIDHT*123]),
			.Valid_Out(CHANNEL124_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL125 (
			.Data_In(Data_In[DATA_WIDHT*125-1:DATA_WIDHT*124]),
			.Kernel0(32'b10111110100100110010100100000111),
			.Kernel1(32'b10111111000101111110010010101011),
			.Kernel2(32'b10111111000100111110101110101010),
			.Kernel3(32'b10111101100011111110010000111111),
			.Kernel4(32'b10111111001000111110001100110110),
			.Kernel5(32'b10111110010010011100101000011111),
			.Kernel6(32'b00111110011000101011100000010001),
			.Kernel7(32'b00111110100100110110111111010001),
			.Kernel8(32'b00111110101001110101100011010011),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*125-1:DATA_WIDHT*124]),
			.Valid_Out(CHANNEL125_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL126 (
			.Data_In(Data_In[DATA_WIDHT*126-1:DATA_WIDHT*125]),
			.Kernel0(32'b10111110100100101110001001011000),
			.Kernel1(32'b10111111000010010010001111000000),
			.Kernel2(32'b10111110111010010001001100111110),
			.Kernel3(32'b10111101110111000110111011110100),
			.Kernel4(32'b10111110010010111001010100101001),
			.Kernel5(32'b00111110000011101101110100000100),
			.Kernel6(32'b00111110111101011101111000111101),
			.Kernel7(32'b00111111000001101010000111000101),
			.Kernel8(32'b00111111000101000110010000001111),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*126-1:DATA_WIDHT*125]),
			.Valid_Out(CHANNEL126_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL127 (
			.Data_In(Data_In[DATA_WIDHT*127-1:DATA_WIDHT*126]),
			.Kernel0(32'b10111111001001000110000011110100),
			.Kernel1(32'b10111111001001101001101101000101),
			.Kernel2(32'b10111111001011101011111000111100),
			.Kernel3(32'b10111101110010100110110100000001),
			.Kernel4(32'b10111110011100001100101110110100),
			.Kernel5(32'b10111110000110100100101000100101),
			.Kernel6(32'b00111101011100111110010010001011),
			.Kernel7(32'b00111110001110000100011110111011),
			.Kernel8(32'b00111111000111100111011101111100),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*127-1:DATA_WIDHT*126]),
			.Valid_Out(CHANNEL127_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL128 (
			.Data_In(Data_In[DATA_WIDHT*128-1:DATA_WIDHT*127]),
			.Kernel0(32'b00111111010011010011011100011000),
			.Kernel1(32'b00111111000011110101100100000000),
			.Kernel2(32'b00111111000000111101111111100110),
			.Kernel3(32'b00111101000011111010011010001001),
			.Kernel4(32'b10111110011000001000000111000110),
			.Kernel5(32'b10111110000001000000100101010011),
			.Kernel6(32'b10111111000000011110011001010000),
			.Kernel7(32'b00111101010010110011101001011100),
			.Kernel8(32'b10111111000010001100001001101101),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*128-1:DATA_WIDHT*127]),
			.Valid_Out(CHANNEL128_Valid_Out)
		);

    
endmodule