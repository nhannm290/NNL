module Convo_Layer6 #(
    parameter DATA_WIDHT = 32,
	parameter IMG_WIDHT = 44,
	parameter IMG_HEIGHT =44
)
(
    input [DATA_WIDHT*64-1:0] Data_In,
    input Valid_In,
    input clk,
    input rst,
    output [DATA_WIDHT*128-1:0] Data_Out,
    output Valid_Out
);
	wire[DATA_WIDHT*64-1:0] Data_Out_Kernel1, Data_Out_Kernel2, Data_Out_Kernel3, Data_Out_Kernel4, Data_Out_Kernel5, Data_Out_Kernel6, Data_Out_Kernel7, Data_Out_Kernel8, Data_Out_Kernel9, Data_Out_Kernel10, Data_Out_Kernel11, Data_Out_Kernel12, Data_Out_Kernel13, Data_Out_Kernel14, Data_Out_Kernel15, Data_Out_Kernel16, Data_Out_Kernel17, Data_Out_Kernel18, Data_Out_Kernel19, Data_Out_Kernel20, Data_Out_Kernel21, Data_Out_Kernel22, Data_Out_Kernel23, Data_Out_Kernel24, Data_Out_Kernel25, Data_Out_Kernel26, Data_Out_Kernel27, Data_Out_Kernel28, Data_Out_Kernel29, Data_Out_Kernel30, Data_Out_Kernel31, Data_Out_Kernel32, Data_Out_Kernel33, Data_Out_Kernel34, Data_Out_Kernel35, Data_Out_Kernel36, Data_Out_Kernel37, Data_Out_Kernel38, Data_Out_Kernel39, Data_Out_Kernel40, Data_Out_Kernel41, Data_Out_Kernel42, Data_Out_Kernel43, Data_Out_Kernel44, Data_Out_Kernel45, Data_Out_Kernel46, Data_Out_Kernel47, Data_Out_Kernel48, Data_Out_Kernel49, Data_Out_Kernel50, Data_Out_Kernel51, Data_Out_Kernel52, Data_Out_Kernel53, Data_Out_Kernel54, Data_Out_Kernel55, Data_Out_Kernel56, Data_Out_Kernel57, Data_Out_Kernel58, Data_Out_Kernel59, Data_Out_Kernel60, Data_Out_Kernel61, Data_Out_Kernel62, Data_Out_Kernel63, Data_Out_Kernel64, Data_Out_Kernel65, Data_Out_Kernel66, Data_Out_Kernel67, Data_Out_Kernel68, Data_Out_Kernel69, Data_Out_Kernel70, Data_Out_Kernel71, Data_Out_Kernel72, Data_Out_Kernel73, Data_Out_Kernel74, Data_Out_Kernel75, Data_Out_Kernel76, Data_Out_Kernel77, Data_Out_Kernel78, Data_Out_Kernel79, Data_Out_Kernel80, Data_Out_Kernel81, Data_Out_Kernel82, Data_Out_Kernel83, Data_Out_Kernel84, Data_Out_Kernel85, Data_Out_Kernel86, Data_Out_Kernel87, Data_Out_Kernel88, Data_Out_Kernel89, Data_Out_Kernel90, Data_Out_Kernel91, Data_Out_Kernel92, Data_Out_Kernel93, Data_Out_Kernel94, Data_Out_Kernel95, Data_Out_Kernel96, Data_Out_Kernel97, Data_Out_Kernel98, Data_Out_Kernel99, Data_Out_Kernel100, Data_Out_Kernel101, Data_Out_Kernel102, Data_Out_Kernel103, Data_Out_Kernel104, Data_Out_Kernel105, Data_Out_Kernel106, Data_Out_Kernel107, Data_Out_Kernel108, Data_Out_Kernel109, Data_Out_Kernel110, Data_Out_Kernel111, Data_Out_Kernel112, Data_Out_Kernel113, Data_Out_Kernel114, Data_Out_Kernel115, Data_Out_Kernel116, Data_Out_Kernel117, Data_Out_Kernel118, Data_Out_Kernel119, Data_Out_Kernel120, Data_Out_Kernel121, Data_Out_Kernel122, Data_Out_Kernel123, Data_Out_Kernel124, Data_Out_Kernel125, Data_Out_Kernel126, Data_Out_Kernel127, Data_Out_Kernel128;
	wire[31:0] add_k1_Data_Out, add_k2_Data_Out, add_k3_Data_Out, add_k4_Data_Out, add_k5_Data_Out, add_k6_Data_Out, add_k7_Data_Out, add_k8_Data_Out, add_k9_Data_Out, add_k10_Data_Out, add_k11_Data_Out, add_k12_Data_Out, add_k13_Data_Out, add_k14_Data_Out, add_k15_Data_Out, add_k16_Data_Out, add_k17_Data_Out, add_k18_Data_Out, add_k19_Data_Out, add_k20_Data_Out, add_k21_Data_Out, add_k22_Data_Out, add_k23_Data_Out, add_k24_Data_Out, add_k25_Data_Out, add_k26_Data_Out, add_k27_Data_Out, add_k28_Data_Out, add_k29_Data_Out, add_k30_Data_Out, add_k31_Data_Out, add_k32_Data_Out, add_k33_Data_Out, add_k34_Data_Out, add_k35_Data_Out, add_k36_Data_Out, add_k37_Data_Out, add_k38_Data_Out, add_k39_Data_Out, add_k40_Data_Out, add_k41_Data_Out, add_k42_Data_Out, add_k43_Data_Out, add_k44_Data_Out, add_k45_Data_Out, add_k46_Data_Out, add_k47_Data_Out, add_k48_Data_Out, add_k49_Data_Out, add_k50_Data_Out, add_k51_Data_Out, add_k52_Data_Out, add_k53_Data_Out, add_k54_Data_Out, add_k55_Data_Out, add_k56_Data_Out, add_k57_Data_Out, add_k58_Data_Out, add_k59_Data_Out, add_k60_Data_Out, add_k61_Data_Out, add_k62_Data_Out, add_k63_Data_Out, add_k64_Data_Out, add_k65_Data_Out, add_k66_Data_Out, add_k67_Data_Out, add_k68_Data_Out, add_k69_Data_Out, add_k70_Data_Out, add_k71_Data_Out, add_k72_Data_Out, add_k73_Data_Out, add_k74_Data_Out, add_k75_Data_Out, add_k76_Data_Out, add_k77_Data_Out, add_k78_Data_Out, add_k79_Data_Out, add_k80_Data_Out, add_k81_Data_Out, add_k82_Data_Out, add_k83_Data_Out, add_k84_Data_Out, add_k85_Data_Out, add_k86_Data_Out, add_k87_Data_Out, add_k88_Data_Out, add_k89_Data_Out, add_k90_Data_Out, add_k91_Data_Out, add_k92_Data_Out, add_k93_Data_Out, add_k94_Data_Out, add_k95_Data_Out, add_k96_Data_Out, add_k97_Data_Out, add_k98_Data_Out, add_k99_Data_Out, add_k100_Data_Out, add_k101_Data_Out, add_k102_Data_Out, add_k103_Data_Out, add_k104_Data_Out, add_k105_Data_Out, add_k106_Data_Out, add_k107_Data_Out, add_k108_Data_Out, add_k109_Data_Out, add_k110_Data_Out, add_k111_Data_Out, add_k112_Data_Out, add_k113_Data_Out, add_k114_Data_Out, add_k115_Data_Out, add_k116_Data_Out, add_k117_Data_Out, add_k118_Data_Out, add_k119_Data_Out, add_k120_Data_Out, add_k121_Data_Out, add_k122_Data_Out, add_k123_Data_Out, add_k124_Data_Out, add_k125_Data_Out, add_k126_Data_Out, add_k127_Data_Out, add_k128_Data_Out;

	wire add_kernel1_Valid_Out, add_kernel2_Valid_Out, add_kernel3_Valid_Out, add_kernel4_Valid_Out, add_kernel5_Valid_Out, add_kernel6_Valid_Out, add_kernel7_Valid_Out, add_kernel8_Valid_Out, add_kernel9_Valid_Out, add_kernel10_Valid_Out, add_kernel11_Valid_Out, add_kernel12_Valid_Out, add_kernel13_Valid_Out, add_kernel14_Valid_Out, add_kernel15_Valid_Out, add_kernel16_Valid_Out, add_kernel17_Valid_Out, add_kernel18_Valid_Out, add_kernel19_Valid_Out, add_kernel20_Valid_Out, add_kernel21_Valid_Out, add_kernel22_Valid_Out, add_kernel23_Valid_Out, add_kernel24_Valid_Out, add_kernel25_Valid_Out, add_kernel26_Valid_Out, add_kernel27_Valid_Out, add_kernel28_Valid_Out, add_kernel29_Valid_Out, add_kernel30_Valid_Out, add_kernel31_Valid_Out, add_kernel32_Valid_Out, add_kernel33_Valid_Out, add_kernel34_Valid_Out, add_kernel35_Valid_Out, add_kernel36_Valid_Out, add_kernel37_Valid_Out, add_kernel38_Valid_Out, add_kernel39_Valid_Out, add_kernel40_Valid_Out, add_kernel41_Valid_Out, add_kernel42_Valid_Out, add_kernel43_Valid_Out, add_kernel44_Valid_Out, add_kernel45_Valid_Out, add_kernel46_Valid_Out, add_kernel47_Valid_Out, add_kernel48_Valid_Out, add_kernel49_Valid_Out, add_kernel50_Valid_Out, add_kernel51_Valid_Out, add_kernel52_Valid_Out, add_kernel53_Valid_Out, add_kernel54_Valid_Out, add_kernel55_Valid_Out, add_kernel56_Valid_Out, add_kernel57_Valid_Out, add_kernel58_Valid_Out, add_kernel59_Valid_Out, add_kernel60_Valid_Out, add_kernel61_Valid_Out, add_kernel62_Valid_Out, add_kernel63_Valid_Out, add_kernel64_Valid_Out, add_kernel65_Valid_Out, add_kernel66_Valid_Out, add_kernel67_Valid_Out, add_kernel68_Valid_Out, add_kernel69_Valid_Out, add_kernel70_Valid_Out, add_kernel71_Valid_Out, add_kernel72_Valid_Out, add_kernel73_Valid_Out, add_kernel74_Valid_Out, add_kernel75_Valid_Out, add_kernel76_Valid_Out, add_kernel77_Valid_Out, add_kernel78_Valid_Out, add_kernel79_Valid_Out, add_kernel80_Valid_Out, add_kernel81_Valid_Out, add_kernel82_Valid_Out, add_kernel83_Valid_Out, add_kernel84_Valid_Out, add_kernel85_Valid_Out, add_kernel86_Valid_Out, add_kernel87_Valid_Out, add_kernel88_Valid_Out, add_kernel89_Valid_Out, add_kernel90_Valid_Out, add_kernel91_Valid_Out, add_kernel92_Valid_Out, add_kernel93_Valid_Out, add_kernel94_Valid_Out, add_kernel95_Valid_Out, add_kernel96_Valid_Out, add_kernel97_Valid_Out, add_kernel98_Valid_Out, add_kernel99_Valid_Out, add_kernel100_Valid_Out, add_kernel101_Valid_Out, add_kernel102_Valid_Out, add_kernel103_Valid_Out, add_kernel104_Valid_Out, add_kernel105_Valid_Out, add_kernel106_Valid_Out, add_kernel107_Valid_Out, add_kernel108_Valid_Out, add_kernel109_Valid_Out, add_kernel110_Valid_Out, add_kernel111_Valid_Out, add_kernel112_Valid_Out, add_kernel113_Valid_Out, add_kernel114_Valid_Out, add_kernel115_Valid_Out, add_kernel116_Valid_Out, add_kernel117_Valid_Out, add_kernel118_Valid_Out, add_kernel119_Valid_Out, add_kernel120_Valid_Out, add_kernel121_Valid_Out, add_kernel122_Valid_Out, add_kernel123_Valid_Out, add_kernel124_Valid_Out, add_kernel125_Valid_Out, add_kernel126_Valid_Out, add_kernel127_Valid_Out, add_kernel128_Valid_Out;

	wire channel1_Kernel1_Valid_Out, channel2_Kernel1_Valid_Out, channel3_Kernel1_Valid_Out, channel4_Kernel1_Valid_Out, channel5_Kernel1_Valid_Out, channel6_Kernel1_Valid_Out, channel7_Kernel1_Valid_Out, channel8_Kernel1_Valid_Out, channel9_Kernel1_Valid_Out, channel10_Kernel1_Valid_Out, channel11_Kernel1_Valid_Out, channel12_Kernel1_Valid_Out, channel13_Kernel1_Valid_Out, channel14_Kernel1_Valid_Out, channel15_Kernel1_Valid_Out, channel16_Kernel1_Valid_Out, channel17_Kernel1_Valid_Out, channel18_Kernel1_Valid_Out, channel19_Kernel1_Valid_Out, channel20_Kernel1_Valid_Out, channel21_Kernel1_Valid_Out, channel22_Kernel1_Valid_Out, channel23_Kernel1_Valid_Out, channel24_Kernel1_Valid_Out, channel25_Kernel1_Valid_Out, channel26_Kernel1_Valid_Out, channel27_Kernel1_Valid_Out, channel28_Kernel1_Valid_Out, channel29_Kernel1_Valid_Out, channel30_Kernel1_Valid_Out, channel31_Kernel1_Valid_Out, channel32_Kernel1_Valid_Out, channel33_Kernel1_Valid_Out, channel34_Kernel1_Valid_Out, channel35_Kernel1_Valid_Out, channel36_Kernel1_Valid_Out, channel37_Kernel1_Valid_Out, channel38_Kernel1_Valid_Out, channel39_Kernel1_Valid_Out, channel40_Kernel1_Valid_Out, channel41_Kernel1_Valid_Out, channel42_Kernel1_Valid_Out, channel43_Kernel1_Valid_Out, channel44_Kernel1_Valid_Out, channel45_Kernel1_Valid_Out, channel46_Kernel1_Valid_Out, channel47_Kernel1_Valid_Out, channel48_Kernel1_Valid_Out, channel49_Kernel1_Valid_Out, channel50_Kernel1_Valid_Out, channel51_Kernel1_Valid_Out, channel52_Kernel1_Valid_Out, channel53_Kernel1_Valid_Out, channel54_Kernel1_Valid_Out, channel55_Kernel1_Valid_Out, channel56_Kernel1_Valid_Out, channel57_Kernel1_Valid_Out, channel58_Kernel1_Valid_Out, channel59_Kernel1_Valid_Out, channel60_Kernel1_Valid_Out, channel61_Kernel1_Valid_Out, channel62_Kernel1_Valid_Out, channel63_Kernel1_Valid_Out, channel64_Kernel1_Valid_Out;

	assign add_kernel1=channel1_Kernel1_Valid_Out & channel2_Kernel1_Valid_Out & channel3_Kernel1_Valid_Out & channel4_Kernel1_Valid_Out & channel5_Kernel1_Valid_Out & channel6_Kernel1_Valid_Out & channel7_Kernel1_Valid_Out & channel8_Kernel1_Valid_Out & channel9_Kernel1_Valid_Out & channel10_Kernel1_Valid_Out & channel11_Kernel1_Valid_Out & channel12_Kernel1_Valid_Out & channel13_Kernel1_Valid_Out & channel14_Kernel1_Valid_Out & channel15_Kernel1_Valid_Out & channel16_Kernel1_Valid_Out & channel17_Kernel1_Valid_Out & channel18_Kernel1_Valid_Out & channel19_Kernel1_Valid_Out & channel20_Kernel1_Valid_Out & channel21_Kernel1_Valid_Out & channel22_Kernel1_Valid_Out & channel23_Kernel1_Valid_Out & channel24_Kernel1_Valid_Out & channel25_Kernel1_Valid_Out & channel26_Kernel1_Valid_Out & channel27_Kernel1_Valid_Out & channel28_Kernel1_Valid_Out & channel29_Kernel1_Valid_Out & channel30_Kernel1_Valid_Out & channel31_Kernel1_Valid_Out & channel32_Kernel1_Valid_Out & channel33_Kernel1_Valid_Out & channel34_Kernel1_Valid_Out & channel35_Kernel1_Valid_Out & channel36_Kernel1_Valid_Out & channel37_Kernel1_Valid_Out & channel38_Kernel1_Valid_Out & channel39_Kernel1_Valid_Out & channel40_Kernel1_Valid_Out & channel41_Kernel1_Valid_Out & channel42_Kernel1_Valid_Out & channel43_Kernel1_Valid_Out & channel44_Kernel1_Valid_Out & channel45_Kernel1_Valid_Out & channel46_Kernel1_Valid_Out & channel47_Kernel1_Valid_Out & channel48_Kernel1_Valid_Out & channel49_Kernel1_Valid_Out & channel50_Kernel1_Valid_Out & channel51_Kernel1_Valid_Out & channel52_Kernel1_Valid_Out & channel53_Kernel1_Valid_Out & channel54_Kernel1_Valid_Out & channel55_Kernel1_Valid_Out & channel56_Kernel1_Valid_Out & channel57_Kernel1_Valid_Out & channel58_Kernel1_Valid_Out & channel59_Kernel1_Valid_Out & channel60_Kernel1_Valid_Out & channel61_Kernel1_Valid_Out & channel62_Kernel1_Valid_Out & channel63_Kernel1_Valid_Out & channel64_Kernel1_Valid_Out;

	wire channel1_Kernel2_Valid_Out, channel2_Kernel2_Valid_Out, channel3_Kernel2_Valid_Out, channel4_Kernel2_Valid_Out, channel5_Kernel2_Valid_Out, channel6_Kernel2_Valid_Out, channel7_Kernel2_Valid_Out, channel8_Kernel2_Valid_Out, channel9_Kernel2_Valid_Out, channel10_Kernel2_Valid_Out, channel11_Kernel2_Valid_Out, channel12_Kernel2_Valid_Out, channel13_Kernel2_Valid_Out, channel14_Kernel2_Valid_Out, channel15_Kernel2_Valid_Out, channel16_Kernel2_Valid_Out, channel17_Kernel2_Valid_Out, channel18_Kernel2_Valid_Out, channel19_Kernel2_Valid_Out, channel20_Kernel2_Valid_Out, channel21_Kernel2_Valid_Out, channel22_Kernel2_Valid_Out, channel23_Kernel2_Valid_Out, channel24_Kernel2_Valid_Out, channel25_Kernel2_Valid_Out, channel26_Kernel2_Valid_Out, channel27_Kernel2_Valid_Out, channel28_Kernel2_Valid_Out, channel29_Kernel2_Valid_Out, channel30_Kernel2_Valid_Out, channel31_Kernel2_Valid_Out, channel32_Kernel2_Valid_Out, channel33_Kernel2_Valid_Out, channel34_Kernel2_Valid_Out, channel35_Kernel2_Valid_Out, channel36_Kernel2_Valid_Out, channel37_Kernel2_Valid_Out, channel38_Kernel2_Valid_Out, channel39_Kernel2_Valid_Out, channel40_Kernel2_Valid_Out, channel41_Kernel2_Valid_Out, channel42_Kernel2_Valid_Out, channel43_Kernel2_Valid_Out, channel44_Kernel2_Valid_Out, channel45_Kernel2_Valid_Out, channel46_Kernel2_Valid_Out, channel47_Kernel2_Valid_Out, channel48_Kernel2_Valid_Out, channel49_Kernel2_Valid_Out, channel50_Kernel2_Valid_Out, channel51_Kernel2_Valid_Out, channel52_Kernel2_Valid_Out, channel53_Kernel2_Valid_Out, channel54_Kernel2_Valid_Out, channel55_Kernel2_Valid_Out, channel56_Kernel2_Valid_Out, channel57_Kernel2_Valid_Out, channel58_Kernel2_Valid_Out, channel59_Kernel2_Valid_Out, channel60_Kernel2_Valid_Out, channel61_Kernel2_Valid_Out, channel62_Kernel2_Valid_Out, channel63_Kernel2_Valid_Out, channel64_Kernel2_Valid_Out;

	assign add_kernel2=channel1_Kernel2_Valid_Out & channel2_Kernel2_Valid_Out & channel3_Kernel2_Valid_Out & channel4_Kernel2_Valid_Out & channel5_Kernel2_Valid_Out & channel6_Kernel2_Valid_Out & channel7_Kernel2_Valid_Out & channel8_Kernel2_Valid_Out & channel9_Kernel2_Valid_Out & channel10_Kernel2_Valid_Out & channel11_Kernel2_Valid_Out & channel12_Kernel2_Valid_Out & channel13_Kernel2_Valid_Out & channel14_Kernel2_Valid_Out & channel15_Kernel2_Valid_Out & channel16_Kernel2_Valid_Out & channel17_Kernel2_Valid_Out & channel18_Kernel2_Valid_Out & channel19_Kernel2_Valid_Out & channel20_Kernel2_Valid_Out & channel21_Kernel2_Valid_Out & channel22_Kernel2_Valid_Out & channel23_Kernel2_Valid_Out & channel24_Kernel2_Valid_Out & channel25_Kernel2_Valid_Out & channel26_Kernel2_Valid_Out & channel27_Kernel2_Valid_Out & channel28_Kernel2_Valid_Out & channel29_Kernel2_Valid_Out & channel30_Kernel2_Valid_Out & channel31_Kernel2_Valid_Out & channel32_Kernel2_Valid_Out & channel33_Kernel2_Valid_Out & channel34_Kernel2_Valid_Out & channel35_Kernel2_Valid_Out & channel36_Kernel2_Valid_Out & channel37_Kernel2_Valid_Out & channel38_Kernel2_Valid_Out & channel39_Kernel2_Valid_Out & channel40_Kernel2_Valid_Out & channel41_Kernel2_Valid_Out & channel42_Kernel2_Valid_Out & channel43_Kernel2_Valid_Out & channel44_Kernel2_Valid_Out & channel45_Kernel2_Valid_Out & channel46_Kernel2_Valid_Out & channel47_Kernel2_Valid_Out & channel48_Kernel2_Valid_Out & channel49_Kernel2_Valid_Out & channel50_Kernel2_Valid_Out & channel51_Kernel2_Valid_Out & channel52_Kernel2_Valid_Out & channel53_Kernel2_Valid_Out & channel54_Kernel2_Valid_Out & channel55_Kernel2_Valid_Out & channel56_Kernel2_Valid_Out & channel57_Kernel2_Valid_Out & channel58_Kernel2_Valid_Out & channel59_Kernel2_Valid_Out & channel60_Kernel2_Valid_Out & channel61_Kernel2_Valid_Out & channel62_Kernel2_Valid_Out & channel63_Kernel2_Valid_Out & channel64_Kernel2_Valid_Out;

	wire channel1_Kernel3_Valid_Out, channel2_Kernel3_Valid_Out, channel3_Kernel3_Valid_Out, channel4_Kernel3_Valid_Out, channel5_Kernel3_Valid_Out, channel6_Kernel3_Valid_Out, channel7_Kernel3_Valid_Out, channel8_Kernel3_Valid_Out, channel9_Kernel3_Valid_Out, channel10_Kernel3_Valid_Out, channel11_Kernel3_Valid_Out, channel12_Kernel3_Valid_Out, channel13_Kernel3_Valid_Out, channel14_Kernel3_Valid_Out, channel15_Kernel3_Valid_Out, channel16_Kernel3_Valid_Out, channel17_Kernel3_Valid_Out, channel18_Kernel3_Valid_Out, channel19_Kernel3_Valid_Out, channel20_Kernel3_Valid_Out, channel21_Kernel3_Valid_Out, channel22_Kernel3_Valid_Out, channel23_Kernel3_Valid_Out, channel24_Kernel3_Valid_Out, channel25_Kernel3_Valid_Out, channel26_Kernel3_Valid_Out, channel27_Kernel3_Valid_Out, channel28_Kernel3_Valid_Out, channel29_Kernel3_Valid_Out, channel30_Kernel3_Valid_Out, channel31_Kernel3_Valid_Out, channel32_Kernel3_Valid_Out, channel33_Kernel3_Valid_Out, channel34_Kernel3_Valid_Out, channel35_Kernel3_Valid_Out, channel36_Kernel3_Valid_Out, channel37_Kernel3_Valid_Out, channel38_Kernel3_Valid_Out, channel39_Kernel3_Valid_Out, channel40_Kernel3_Valid_Out, channel41_Kernel3_Valid_Out, channel42_Kernel3_Valid_Out, channel43_Kernel3_Valid_Out, channel44_Kernel3_Valid_Out, channel45_Kernel3_Valid_Out, channel46_Kernel3_Valid_Out, channel47_Kernel3_Valid_Out, channel48_Kernel3_Valid_Out, channel49_Kernel3_Valid_Out, channel50_Kernel3_Valid_Out, channel51_Kernel3_Valid_Out, channel52_Kernel3_Valid_Out, channel53_Kernel3_Valid_Out, channel54_Kernel3_Valid_Out, channel55_Kernel3_Valid_Out, channel56_Kernel3_Valid_Out, channel57_Kernel3_Valid_Out, channel58_Kernel3_Valid_Out, channel59_Kernel3_Valid_Out, channel60_Kernel3_Valid_Out, channel61_Kernel3_Valid_Out, channel62_Kernel3_Valid_Out, channel63_Kernel3_Valid_Out, channel64_Kernel3_Valid_Out;

	assign add_kernel3=channel1_Kernel3_Valid_Out & channel2_Kernel3_Valid_Out & channel3_Kernel3_Valid_Out & channel4_Kernel3_Valid_Out & channel5_Kernel3_Valid_Out & channel6_Kernel3_Valid_Out & channel7_Kernel3_Valid_Out & channel8_Kernel3_Valid_Out & channel9_Kernel3_Valid_Out & channel10_Kernel3_Valid_Out & channel11_Kernel3_Valid_Out & channel12_Kernel3_Valid_Out & channel13_Kernel3_Valid_Out & channel14_Kernel3_Valid_Out & channel15_Kernel3_Valid_Out & channel16_Kernel3_Valid_Out & channel17_Kernel3_Valid_Out & channel18_Kernel3_Valid_Out & channel19_Kernel3_Valid_Out & channel20_Kernel3_Valid_Out & channel21_Kernel3_Valid_Out & channel22_Kernel3_Valid_Out & channel23_Kernel3_Valid_Out & channel24_Kernel3_Valid_Out & channel25_Kernel3_Valid_Out & channel26_Kernel3_Valid_Out & channel27_Kernel3_Valid_Out & channel28_Kernel3_Valid_Out & channel29_Kernel3_Valid_Out & channel30_Kernel3_Valid_Out & channel31_Kernel3_Valid_Out & channel32_Kernel3_Valid_Out & channel33_Kernel3_Valid_Out & channel34_Kernel3_Valid_Out & channel35_Kernel3_Valid_Out & channel36_Kernel3_Valid_Out & channel37_Kernel3_Valid_Out & channel38_Kernel3_Valid_Out & channel39_Kernel3_Valid_Out & channel40_Kernel3_Valid_Out & channel41_Kernel3_Valid_Out & channel42_Kernel3_Valid_Out & channel43_Kernel3_Valid_Out & channel44_Kernel3_Valid_Out & channel45_Kernel3_Valid_Out & channel46_Kernel3_Valid_Out & channel47_Kernel3_Valid_Out & channel48_Kernel3_Valid_Out & channel49_Kernel3_Valid_Out & channel50_Kernel3_Valid_Out & channel51_Kernel3_Valid_Out & channel52_Kernel3_Valid_Out & channel53_Kernel3_Valid_Out & channel54_Kernel3_Valid_Out & channel55_Kernel3_Valid_Out & channel56_Kernel3_Valid_Out & channel57_Kernel3_Valid_Out & channel58_Kernel3_Valid_Out & channel59_Kernel3_Valid_Out & channel60_Kernel3_Valid_Out & channel61_Kernel3_Valid_Out & channel62_Kernel3_Valid_Out & channel63_Kernel3_Valid_Out & channel64_Kernel3_Valid_Out;

	wire channel1_Kernel4_Valid_Out, channel2_Kernel4_Valid_Out, channel3_Kernel4_Valid_Out, channel4_Kernel4_Valid_Out, channel5_Kernel4_Valid_Out, channel6_Kernel4_Valid_Out, channel7_Kernel4_Valid_Out, channel8_Kernel4_Valid_Out, channel9_Kernel4_Valid_Out, channel10_Kernel4_Valid_Out, channel11_Kernel4_Valid_Out, channel12_Kernel4_Valid_Out, channel13_Kernel4_Valid_Out, channel14_Kernel4_Valid_Out, channel15_Kernel4_Valid_Out, channel16_Kernel4_Valid_Out, channel17_Kernel4_Valid_Out, channel18_Kernel4_Valid_Out, channel19_Kernel4_Valid_Out, channel20_Kernel4_Valid_Out, channel21_Kernel4_Valid_Out, channel22_Kernel4_Valid_Out, channel23_Kernel4_Valid_Out, channel24_Kernel4_Valid_Out, channel25_Kernel4_Valid_Out, channel26_Kernel4_Valid_Out, channel27_Kernel4_Valid_Out, channel28_Kernel4_Valid_Out, channel29_Kernel4_Valid_Out, channel30_Kernel4_Valid_Out, channel31_Kernel4_Valid_Out, channel32_Kernel4_Valid_Out, channel33_Kernel4_Valid_Out, channel34_Kernel4_Valid_Out, channel35_Kernel4_Valid_Out, channel36_Kernel4_Valid_Out, channel37_Kernel4_Valid_Out, channel38_Kernel4_Valid_Out, channel39_Kernel4_Valid_Out, channel40_Kernel4_Valid_Out, channel41_Kernel4_Valid_Out, channel42_Kernel4_Valid_Out, channel43_Kernel4_Valid_Out, channel44_Kernel4_Valid_Out, channel45_Kernel4_Valid_Out, channel46_Kernel4_Valid_Out, channel47_Kernel4_Valid_Out, channel48_Kernel4_Valid_Out, channel49_Kernel4_Valid_Out, channel50_Kernel4_Valid_Out, channel51_Kernel4_Valid_Out, channel52_Kernel4_Valid_Out, channel53_Kernel4_Valid_Out, channel54_Kernel4_Valid_Out, channel55_Kernel4_Valid_Out, channel56_Kernel4_Valid_Out, channel57_Kernel4_Valid_Out, channel58_Kernel4_Valid_Out, channel59_Kernel4_Valid_Out, channel60_Kernel4_Valid_Out, channel61_Kernel4_Valid_Out, channel62_Kernel4_Valid_Out, channel63_Kernel4_Valid_Out, channel64_Kernel4_Valid_Out;

	assign add_kernel4=channel1_Kernel4_Valid_Out & channel2_Kernel4_Valid_Out & channel3_Kernel4_Valid_Out & channel4_Kernel4_Valid_Out & channel5_Kernel4_Valid_Out & channel6_Kernel4_Valid_Out & channel7_Kernel4_Valid_Out & channel8_Kernel4_Valid_Out & channel9_Kernel4_Valid_Out & channel10_Kernel4_Valid_Out & channel11_Kernel4_Valid_Out & channel12_Kernel4_Valid_Out & channel13_Kernel4_Valid_Out & channel14_Kernel4_Valid_Out & channel15_Kernel4_Valid_Out & channel16_Kernel4_Valid_Out & channel17_Kernel4_Valid_Out & channel18_Kernel4_Valid_Out & channel19_Kernel4_Valid_Out & channel20_Kernel4_Valid_Out & channel21_Kernel4_Valid_Out & channel22_Kernel4_Valid_Out & channel23_Kernel4_Valid_Out & channel24_Kernel4_Valid_Out & channel25_Kernel4_Valid_Out & channel26_Kernel4_Valid_Out & channel27_Kernel4_Valid_Out & channel28_Kernel4_Valid_Out & channel29_Kernel4_Valid_Out & channel30_Kernel4_Valid_Out & channel31_Kernel4_Valid_Out & channel32_Kernel4_Valid_Out & channel33_Kernel4_Valid_Out & channel34_Kernel4_Valid_Out & channel35_Kernel4_Valid_Out & channel36_Kernel4_Valid_Out & channel37_Kernel4_Valid_Out & channel38_Kernel4_Valid_Out & channel39_Kernel4_Valid_Out & channel40_Kernel4_Valid_Out & channel41_Kernel4_Valid_Out & channel42_Kernel4_Valid_Out & channel43_Kernel4_Valid_Out & channel44_Kernel4_Valid_Out & channel45_Kernel4_Valid_Out & channel46_Kernel4_Valid_Out & channel47_Kernel4_Valid_Out & channel48_Kernel4_Valid_Out & channel49_Kernel4_Valid_Out & channel50_Kernel4_Valid_Out & channel51_Kernel4_Valid_Out & channel52_Kernel4_Valid_Out & channel53_Kernel4_Valid_Out & channel54_Kernel4_Valid_Out & channel55_Kernel4_Valid_Out & channel56_Kernel4_Valid_Out & channel57_Kernel4_Valid_Out & channel58_Kernel4_Valid_Out & channel59_Kernel4_Valid_Out & channel60_Kernel4_Valid_Out & channel61_Kernel4_Valid_Out & channel62_Kernel4_Valid_Out & channel63_Kernel4_Valid_Out & channel64_Kernel4_Valid_Out;

	wire channel1_Kernel5_Valid_Out, channel2_Kernel5_Valid_Out, channel3_Kernel5_Valid_Out, channel4_Kernel5_Valid_Out, channel5_Kernel5_Valid_Out, channel6_Kernel5_Valid_Out, channel7_Kernel5_Valid_Out, channel8_Kernel5_Valid_Out, channel9_Kernel5_Valid_Out, channel10_Kernel5_Valid_Out, channel11_Kernel5_Valid_Out, channel12_Kernel5_Valid_Out, channel13_Kernel5_Valid_Out, channel14_Kernel5_Valid_Out, channel15_Kernel5_Valid_Out, channel16_Kernel5_Valid_Out, channel17_Kernel5_Valid_Out, channel18_Kernel5_Valid_Out, channel19_Kernel5_Valid_Out, channel20_Kernel5_Valid_Out, channel21_Kernel5_Valid_Out, channel22_Kernel5_Valid_Out, channel23_Kernel5_Valid_Out, channel24_Kernel5_Valid_Out, channel25_Kernel5_Valid_Out, channel26_Kernel5_Valid_Out, channel27_Kernel5_Valid_Out, channel28_Kernel5_Valid_Out, channel29_Kernel5_Valid_Out, channel30_Kernel5_Valid_Out, channel31_Kernel5_Valid_Out, channel32_Kernel5_Valid_Out, channel33_Kernel5_Valid_Out, channel34_Kernel5_Valid_Out, channel35_Kernel5_Valid_Out, channel36_Kernel5_Valid_Out, channel37_Kernel5_Valid_Out, channel38_Kernel5_Valid_Out, channel39_Kernel5_Valid_Out, channel40_Kernel5_Valid_Out, channel41_Kernel5_Valid_Out, channel42_Kernel5_Valid_Out, channel43_Kernel5_Valid_Out, channel44_Kernel5_Valid_Out, channel45_Kernel5_Valid_Out, channel46_Kernel5_Valid_Out, channel47_Kernel5_Valid_Out, channel48_Kernel5_Valid_Out, channel49_Kernel5_Valid_Out, channel50_Kernel5_Valid_Out, channel51_Kernel5_Valid_Out, channel52_Kernel5_Valid_Out, channel53_Kernel5_Valid_Out, channel54_Kernel5_Valid_Out, channel55_Kernel5_Valid_Out, channel56_Kernel5_Valid_Out, channel57_Kernel5_Valid_Out, channel58_Kernel5_Valid_Out, channel59_Kernel5_Valid_Out, channel60_Kernel5_Valid_Out, channel61_Kernel5_Valid_Out, channel62_Kernel5_Valid_Out, channel63_Kernel5_Valid_Out, channel64_Kernel5_Valid_Out;

	assign add_kernel5=channel1_Kernel5_Valid_Out & channel2_Kernel5_Valid_Out & channel3_Kernel5_Valid_Out & channel4_Kernel5_Valid_Out & channel5_Kernel5_Valid_Out & channel6_Kernel5_Valid_Out & channel7_Kernel5_Valid_Out & channel8_Kernel5_Valid_Out & channel9_Kernel5_Valid_Out & channel10_Kernel5_Valid_Out & channel11_Kernel5_Valid_Out & channel12_Kernel5_Valid_Out & channel13_Kernel5_Valid_Out & channel14_Kernel5_Valid_Out & channel15_Kernel5_Valid_Out & channel16_Kernel5_Valid_Out & channel17_Kernel5_Valid_Out & channel18_Kernel5_Valid_Out & channel19_Kernel5_Valid_Out & channel20_Kernel5_Valid_Out & channel21_Kernel5_Valid_Out & channel22_Kernel5_Valid_Out & channel23_Kernel5_Valid_Out & channel24_Kernel5_Valid_Out & channel25_Kernel5_Valid_Out & channel26_Kernel5_Valid_Out & channel27_Kernel5_Valid_Out & channel28_Kernel5_Valid_Out & channel29_Kernel5_Valid_Out & channel30_Kernel5_Valid_Out & channel31_Kernel5_Valid_Out & channel32_Kernel5_Valid_Out & channel33_Kernel5_Valid_Out & channel34_Kernel5_Valid_Out & channel35_Kernel5_Valid_Out & channel36_Kernel5_Valid_Out & channel37_Kernel5_Valid_Out & channel38_Kernel5_Valid_Out & channel39_Kernel5_Valid_Out & channel40_Kernel5_Valid_Out & channel41_Kernel5_Valid_Out & channel42_Kernel5_Valid_Out & channel43_Kernel5_Valid_Out & channel44_Kernel5_Valid_Out & channel45_Kernel5_Valid_Out & channel46_Kernel5_Valid_Out & channel47_Kernel5_Valid_Out & channel48_Kernel5_Valid_Out & channel49_Kernel5_Valid_Out & channel50_Kernel5_Valid_Out & channel51_Kernel5_Valid_Out & channel52_Kernel5_Valid_Out & channel53_Kernel5_Valid_Out & channel54_Kernel5_Valid_Out & channel55_Kernel5_Valid_Out & channel56_Kernel5_Valid_Out & channel57_Kernel5_Valid_Out & channel58_Kernel5_Valid_Out & channel59_Kernel5_Valid_Out & channel60_Kernel5_Valid_Out & channel61_Kernel5_Valid_Out & channel62_Kernel5_Valid_Out & channel63_Kernel5_Valid_Out & channel64_Kernel5_Valid_Out;

	wire channel1_Kernel6_Valid_Out, channel2_Kernel6_Valid_Out, channel3_Kernel6_Valid_Out, channel4_Kernel6_Valid_Out, channel5_Kernel6_Valid_Out, channel6_Kernel6_Valid_Out, channel7_Kernel6_Valid_Out, channel8_Kernel6_Valid_Out, channel9_Kernel6_Valid_Out, channel10_Kernel6_Valid_Out, channel11_Kernel6_Valid_Out, channel12_Kernel6_Valid_Out, channel13_Kernel6_Valid_Out, channel14_Kernel6_Valid_Out, channel15_Kernel6_Valid_Out, channel16_Kernel6_Valid_Out, channel17_Kernel6_Valid_Out, channel18_Kernel6_Valid_Out, channel19_Kernel6_Valid_Out, channel20_Kernel6_Valid_Out, channel21_Kernel6_Valid_Out, channel22_Kernel6_Valid_Out, channel23_Kernel6_Valid_Out, channel24_Kernel6_Valid_Out, channel25_Kernel6_Valid_Out, channel26_Kernel6_Valid_Out, channel27_Kernel6_Valid_Out, channel28_Kernel6_Valid_Out, channel29_Kernel6_Valid_Out, channel30_Kernel6_Valid_Out, channel31_Kernel6_Valid_Out, channel32_Kernel6_Valid_Out, channel33_Kernel6_Valid_Out, channel34_Kernel6_Valid_Out, channel35_Kernel6_Valid_Out, channel36_Kernel6_Valid_Out, channel37_Kernel6_Valid_Out, channel38_Kernel6_Valid_Out, channel39_Kernel6_Valid_Out, channel40_Kernel6_Valid_Out, channel41_Kernel6_Valid_Out, channel42_Kernel6_Valid_Out, channel43_Kernel6_Valid_Out, channel44_Kernel6_Valid_Out, channel45_Kernel6_Valid_Out, channel46_Kernel6_Valid_Out, channel47_Kernel6_Valid_Out, channel48_Kernel6_Valid_Out, channel49_Kernel6_Valid_Out, channel50_Kernel6_Valid_Out, channel51_Kernel6_Valid_Out, channel52_Kernel6_Valid_Out, channel53_Kernel6_Valid_Out, channel54_Kernel6_Valid_Out, channel55_Kernel6_Valid_Out, channel56_Kernel6_Valid_Out, channel57_Kernel6_Valid_Out, channel58_Kernel6_Valid_Out, channel59_Kernel6_Valid_Out, channel60_Kernel6_Valid_Out, channel61_Kernel6_Valid_Out, channel62_Kernel6_Valid_Out, channel63_Kernel6_Valid_Out, channel64_Kernel6_Valid_Out;

	assign add_kernel6=channel1_Kernel6_Valid_Out & channel2_Kernel6_Valid_Out & channel3_Kernel6_Valid_Out & channel4_Kernel6_Valid_Out & channel5_Kernel6_Valid_Out & channel6_Kernel6_Valid_Out & channel7_Kernel6_Valid_Out & channel8_Kernel6_Valid_Out & channel9_Kernel6_Valid_Out & channel10_Kernel6_Valid_Out & channel11_Kernel6_Valid_Out & channel12_Kernel6_Valid_Out & channel13_Kernel6_Valid_Out & channel14_Kernel6_Valid_Out & channel15_Kernel6_Valid_Out & channel16_Kernel6_Valid_Out & channel17_Kernel6_Valid_Out & channel18_Kernel6_Valid_Out & channel19_Kernel6_Valid_Out & channel20_Kernel6_Valid_Out & channel21_Kernel6_Valid_Out & channel22_Kernel6_Valid_Out & channel23_Kernel6_Valid_Out & channel24_Kernel6_Valid_Out & channel25_Kernel6_Valid_Out & channel26_Kernel6_Valid_Out & channel27_Kernel6_Valid_Out & channel28_Kernel6_Valid_Out & channel29_Kernel6_Valid_Out & channel30_Kernel6_Valid_Out & channel31_Kernel6_Valid_Out & channel32_Kernel6_Valid_Out & channel33_Kernel6_Valid_Out & channel34_Kernel6_Valid_Out & channel35_Kernel6_Valid_Out & channel36_Kernel6_Valid_Out & channel37_Kernel6_Valid_Out & channel38_Kernel6_Valid_Out & channel39_Kernel6_Valid_Out & channel40_Kernel6_Valid_Out & channel41_Kernel6_Valid_Out & channel42_Kernel6_Valid_Out & channel43_Kernel6_Valid_Out & channel44_Kernel6_Valid_Out & channel45_Kernel6_Valid_Out & channel46_Kernel6_Valid_Out & channel47_Kernel6_Valid_Out & channel48_Kernel6_Valid_Out & channel49_Kernel6_Valid_Out & channel50_Kernel6_Valid_Out & channel51_Kernel6_Valid_Out & channel52_Kernel6_Valid_Out & channel53_Kernel6_Valid_Out & channel54_Kernel6_Valid_Out & channel55_Kernel6_Valid_Out & channel56_Kernel6_Valid_Out & channel57_Kernel6_Valid_Out & channel58_Kernel6_Valid_Out & channel59_Kernel6_Valid_Out & channel60_Kernel6_Valid_Out & channel61_Kernel6_Valid_Out & channel62_Kernel6_Valid_Out & channel63_Kernel6_Valid_Out & channel64_Kernel6_Valid_Out;

	wire channel1_Kernel7_Valid_Out, channel2_Kernel7_Valid_Out, channel3_Kernel7_Valid_Out, channel4_Kernel7_Valid_Out, channel5_Kernel7_Valid_Out, channel6_Kernel7_Valid_Out, channel7_Kernel7_Valid_Out, channel8_Kernel7_Valid_Out, channel9_Kernel7_Valid_Out, channel10_Kernel7_Valid_Out, channel11_Kernel7_Valid_Out, channel12_Kernel7_Valid_Out, channel13_Kernel7_Valid_Out, channel14_Kernel7_Valid_Out, channel15_Kernel7_Valid_Out, channel16_Kernel7_Valid_Out, channel17_Kernel7_Valid_Out, channel18_Kernel7_Valid_Out, channel19_Kernel7_Valid_Out, channel20_Kernel7_Valid_Out, channel21_Kernel7_Valid_Out, channel22_Kernel7_Valid_Out, channel23_Kernel7_Valid_Out, channel24_Kernel7_Valid_Out, channel25_Kernel7_Valid_Out, channel26_Kernel7_Valid_Out, channel27_Kernel7_Valid_Out, channel28_Kernel7_Valid_Out, channel29_Kernel7_Valid_Out, channel30_Kernel7_Valid_Out, channel31_Kernel7_Valid_Out, channel32_Kernel7_Valid_Out, channel33_Kernel7_Valid_Out, channel34_Kernel7_Valid_Out, channel35_Kernel7_Valid_Out, channel36_Kernel7_Valid_Out, channel37_Kernel7_Valid_Out, channel38_Kernel7_Valid_Out, channel39_Kernel7_Valid_Out, channel40_Kernel7_Valid_Out, channel41_Kernel7_Valid_Out, channel42_Kernel7_Valid_Out, channel43_Kernel7_Valid_Out, channel44_Kernel7_Valid_Out, channel45_Kernel7_Valid_Out, channel46_Kernel7_Valid_Out, channel47_Kernel7_Valid_Out, channel48_Kernel7_Valid_Out, channel49_Kernel7_Valid_Out, channel50_Kernel7_Valid_Out, channel51_Kernel7_Valid_Out, channel52_Kernel7_Valid_Out, channel53_Kernel7_Valid_Out, channel54_Kernel7_Valid_Out, channel55_Kernel7_Valid_Out, channel56_Kernel7_Valid_Out, channel57_Kernel7_Valid_Out, channel58_Kernel7_Valid_Out, channel59_Kernel7_Valid_Out, channel60_Kernel7_Valid_Out, channel61_Kernel7_Valid_Out, channel62_Kernel7_Valid_Out, channel63_Kernel7_Valid_Out, channel64_Kernel7_Valid_Out;

	assign add_kernel7=channel1_Kernel7_Valid_Out & channel2_Kernel7_Valid_Out & channel3_Kernel7_Valid_Out & channel4_Kernel7_Valid_Out & channel5_Kernel7_Valid_Out & channel6_Kernel7_Valid_Out & channel7_Kernel7_Valid_Out & channel8_Kernel7_Valid_Out & channel9_Kernel7_Valid_Out & channel10_Kernel7_Valid_Out & channel11_Kernel7_Valid_Out & channel12_Kernel7_Valid_Out & channel13_Kernel7_Valid_Out & channel14_Kernel7_Valid_Out & channel15_Kernel7_Valid_Out & channel16_Kernel7_Valid_Out & channel17_Kernel7_Valid_Out & channel18_Kernel7_Valid_Out & channel19_Kernel7_Valid_Out & channel20_Kernel7_Valid_Out & channel21_Kernel7_Valid_Out & channel22_Kernel7_Valid_Out & channel23_Kernel7_Valid_Out & channel24_Kernel7_Valid_Out & channel25_Kernel7_Valid_Out & channel26_Kernel7_Valid_Out & channel27_Kernel7_Valid_Out & channel28_Kernel7_Valid_Out & channel29_Kernel7_Valid_Out & channel30_Kernel7_Valid_Out & channel31_Kernel7_Valid_Out & channel32_Kernel7_Valid_Out & channel33_Kernel7_Valid_Out & channel34_Kernel7_Valid_Out & channel35_Kernel7_Valid_Out & channel36_Kernel7_Valid_Out & channel37_Kernel7_Valid_Out & channel38_Kernel7_Valid_Out & channel39_Kernel7_Valid_Out & channel40_Kernel7_Valid_Out & channel41_Kernel7_Valid_Out & channel42_Kernel7_Valid_Out & channel43_Kernel7_Valid_Out & channel44_Kernel7_Valid_Out & channel45_Kernel7_Valid_Out & channel46_Kernel7_Valid_Out & channel47_Kernel7_Valid_Out & channel48_Kernel7_Valid_Out & channel49_Kernel7_Valid_Out & channel50_Kernel7_Valid_Out & channel51_Kernel7_Valid_Out & channel52_Kernel7_Valid_Out & channel53_Kernel7_Valid_Out & channel54_Kernel7_Valid_Out & channel55_Kernel7_Valid_Out & channel56_Kernel7_Valid_Out & channel57_Kernel7_Valid_Out & channel58_Kernel7_Valid_Out & channel59_Kernel7_Valid_Out & channel60_Kernel7_Valid_Out & channel61_Kernel7_Valid_Out & channel62_Kernel7_Valid_Out & channel63_Kernel7_Valid_Out & channel64_Kernel7_Valid_Out;

	wire channel1_Kernel8_Valid_Out, channel2_Kernel8_Valid_Out, channel3_Kernel8_Valid_Out, channel4_Kernel8_Valid_Out, channel5_Kernel8_Valid_Out, channel6_Kernel8_Valid_Out, channel7_Kernel8_Valid_Out, channel8_Kernel8_Valid_Out, channel9_Kernel8_Valid_Out, channel10_Kernel8_Valid_Out, channel11_Kernel8_Valid_Out, channel12_Kernel8_Valid_Out, channel13_Kernel8_Valid_Out, channel14_Kernel8_Valid_Out, channel15_Kernel8_Valid_Out, channel16_Kernel8_Valid_Out, channel17_Kernel8_Valid_Out, channel18_Kernel8_Valid_Out, channel19_Kernel8_Valid_Out, channel20_Kernel8_Valid_Out, channel21_Kernel8_Valid_Out, channel22_Kernel8_Valid_Out, channel23_Kernel8_Valid_Out, channel24_Kernel8_Valid_Out, channel25_Kernel8_Valid_Out, channel26_Kernel8_Valid_Out, channel27_Kernel8_Valid_Out, channel28_Kernel8_Valid_Out, channel29_Kernel8_Valid_Out, channel30_Kernel8_Valid_Out, channel31_Kernel8_Valid_Out, channel32_Kernel8_Valid_Out, channel33_Kernel8_Valid_Out, channel34_Kernel8_Valid_Out, channel35_Kernel8_Valid_Out, channel36_Kernel8_Valid_Out, channel37_Kernel8_Valid_Out, channel38_Kernel8_Valid_Out, channel39_Kernel8_Valid_Out, channel40_Kernel8_Valid_Out, channel41_Kernel8_Valid_Out, channel42_Kernel8_Valid_Out, channel43_Kernel8_Valid_Out, channel44_Kernel8_Valid_Out, channel45_Kernel8_Valid_Out, channel46_Kernel8_Valid_Out, channel47_Kernel8_Valid_Out, channel48_Kernel8_Valid_Out, channel49_Kernel8_Valid_Out, channel50_Kernel8_Valid_Out, channel51_Kernel8_Valid_Out, channel52_Kernel8_Valid_Out, channel53_Kernel8_Valid_Out, channel54_Kernel8_Valid_Out, channel55_Kernel8_Valid_Out, channel56_Kernel8_Valid_Out, channel57_Kernel8_Valid_Out, channel58_Kernel8_Valid_Out, channel59_Kernel8_Valid_Out, channel60_Kernel8_Valid_Out, channel61_Kernel8_Valid_Out, channel62_Kernel8_Valid_Out, channel63_Kernel8_Valid_Out, channel64_Kernel8_Valid_Out;

	assign add_kernel8=channel1_Kernel8_Valid_Out & channel2_Kernel8_Valid_Out & channel3_Kernel8_Valid_Out & channel4_Kernel8_Valid_Out & channel5_Kernel8_Valid_Out & channel6_Kernel8_Valid_Out & channel7_Kernel8_Valid_Out & channel8_Kernel8_Valid_Out & channel9_Kernel8_Valid_Out & channel10_Kernel8_Valid_Out & channel11_Kernel8_Valid_Out & channel12_Kernel8_Valid_Out & channel13_Kernel8_Valid_Out & channel14_Kernel8_Valid_Out & channel15_Kernel8_Valid_Out & channel16_Kernel8_Valid_Out & channel17_Kernel8_Valid_Out & channel18_Kernel8_Valid_Out & channel19_Kernel8_Valid_Out & channel20_Kernel8_Valid_Out & channel21_Kernel8_Valid_Out & channel22_Kernel8_Valid_Out & channel23_Kernel8_Valid_Out & channel24_Kernel8_Valid_Out & channel25_Kernel8_Valid_Out & channel26_Kernel8_Valid_Out & channel27_Kernel8_Valid_Out & channel28_Kernel8_Valid_Out & channel29_Kernel8_Valid_Out & channel30_Kernel8_Valid_Out & channel31_Kernel8_Valid_Out & channel32_Kernel8_Valid_Out & channel33_Kernel8_Valid_Out & channel34_Kernel8_Valid_Out & channel35_Kernel8_Valid_Out & channel36_Kernel8_Valid_Out & channel37_Kernel8_Valid_Out & channel38_Kernel8_Valid_Out & channel39_Kernel8_Valid_Out & channel40_Kernel8_Valid_Out & channel41_Kernel8_Valid_Out & channel42_Kernel8_Valid_Out & channel43_Kernel8_Valid_Out & channel44_Kernel8_Valid_Out & channel45_Kernel8_Valid_Out & channel46_Kernel8_Valid_Out & channel47_Kernel8_Valid_Out & channel48_Kernel8_Valid_Out & channel49_Kernel8_Valid_Out & channel50_Kernel8_Valid_Out & channel51_Kernel8_Valid_Out & channel52_Kernel8_Valid_Out & channel53_Kernel8_Valid_Out & channel54_Kernel8_Valid_Out & channel55_Kernel8_Valid_Out & channel56_Kernel8_Valid_Out & channel57_Kernel8_Valid_Out & channel58_Kernel8_Valid_Out & channel59_Kernel8_Valid_Out & channel60_Kernel8_Valid_Out & channel61_Kernel8_Valid_Out & channel62_Kernel8_Valid_Out & channel63_Kernel8_Valid_Out & channel64_Kernel8_Valid_Out;

	wire channel1_Kernel9_Valid_Out, channel2_Kernel9_Valid_Out, channel3_Kernel9_Valid_Out, channel4_Kernel9_Valid_Out, channel5_Kernel9_Valid_Out, channel6_Kernel9_Valid_Out, channel7_Kernel9_Valid_Out, channel8_Kernel9_Valid_Out, channel9_Kernel9_Valid_Out, channel10_Kernel9_Valid_Out, channel11_Kernel9_Valid_Out, channel12_Kernel9_Valid_Out, channel13_Kernel9_Valid_Out, channel14_Kernel9_Valid_Out, channel15_Kernel9_Valid_Out, channel16_Kernel9_Valid_Out, channel17_Kernel9_Valid_Out, channel18_Kernel9_Valid_Out, channel19_Kernel9_Valid_Out, channel20_Kernel9_Valid_Out, channel21_Kernel9_Valid_Out, channel22_Kernel9_Valid_Out, channel23_Kernel9_Valid_Out, channel24_Kernel9_Valid_Out, channel25_Kernel9_Valid_Out, channel26_Kernel9_Valid_Out, channel27_Kernel9_Valid_Out, channel28_Kernel9_Valid_Out, channel29_Kernel9_Valid_Out, channel30_Kernel9_Valid_Out, channel31_Kernel9_Valid_Out, channel32_Kernel9_Valid_Out, channel33_Kernel9_Valid_Out, channel34_Kernel9_Valid_Out, channel35_Kernel9_Valid_Out, channel36_Kernel9_Valid_Out, channel37_Kernel9_Valid_Out, channel38_Kernel9_Valid_Out, channel39_Kernel9_Valid_Out, channel40_Kernel9_Valid_Out, channel41_Kernel9_Valid_Out, channel42_Kernel9_Valid_Out, channel43_Kernel9_Valid_Out, channel44_Kernel9_Valid_Out, channel45_Kernel9_Valid_Out, channel46_Kernel9_Valid_Out, channel47_Kernel9_Valid_Out, channel48_Kernel9_Valid_Out, channel49_Kernel9_Valid_Out, channel50_Kernel9_Valid_Out, channel51_Kernel9_Valid_Out, channel52_Kernel9_Valid_Out, channel53_Kernel9_Valid_Out, channel54_Kernel9_Valid_Out, channel55_Kernel9_Valid_Out, channel56_Kernel9_Valid_Out, channel57_Kernel9_Valid_Out, channel58_Kernel9_Valid_Out, channel59_Kernel9_Valid_Out, channel60_Kernel9_Valid_Out, channel61_Kernel9_Valid_Out, channel62_Kernel9_Valid_Out, channel63_Kernel9_Valid_Out, channel64_Kernel9_Valid_Out;

	assign add_kernel9=channel1_Kernel9_Valid_Out & channel2_Kernel9_Valid_Out & channel3_Kernel9_Valid_Out & channel4_Kernel9_Valid_Out & channel5_Kernel9_Valid_Out & channel6_Kernel9_Valid_Out & channel7_Kernel9_Valid_Out & channel8_Kernel9_Valid_Out & channel9_Kernel9_Valid_Out & channel10_Kernel9_Valid_Out & channel11_Kernel9_Valid_Out & channel12_Kernel9_Valid_Out & channel13_Kernel9_Valid_Out & channel14_Kernel9_Valid_Out & channel15_Kernel9_Valid_Out & channel16_Kernel9_Valid_Out & channel17_Kernel9_Valid_Out & channel18_Kernel9_Valid_Out & channel19_Kernel9_Valid_Out & channel20_Kernel9_Valid_Out & channel21_Kernel9_Valid_Out & channel22_Kernel9_Valid_Out & channel23_Kernel9_Valid_Out & channel24_Kernel9_Valid_Out & channel25_Kernel9_Valid_Out & channel26_Kernel9_Valid_Out & channel27_Kernel9_Valid_Out & channel28_Kernel9_Valid_Out & channel29_Kernel9_Valid_Out & channel30_Kernel9_Valid_Out & channel31_Kernel9_Valid_Out & channel32_Kernel9_Valid_Out & channel33_Kernel9_Valid_Out & channel34_Kernel9_Valid_Out & channel35_Kernel9_Valid_Out & channel36_Kernel9_Valid_Out & channel37_Kernel9_Valid_Out & channel38_Kernel9_Valid_Out & channel39_Kernel9_Valid_Out & channel40_Kernel9_Valid_Out & channel41_Kernel9_Valid_Out & channel42_Kernel9_Valid_Out & channel43_Kernel9_Valid_Out & channel44_Kernel9_Valid_Out & channel45_Kernel9_Valid_Out & channel46_Kernel9_Valid_Out & channel47_Kernel9_Valid_Out & channel48_Kernel9_Valid_Out & channel49_Kernel9_Valid_Out & channel50_Kernel9_Valid_Out & channel51_Kernel9_Valid_Out & channel52_Kernel9_Valid_Out & channel53_Kernel9_Valid_Out & channel54_Kernel9_Valid_Out & channel55_Kernel9_Valid_Out & channel56_Kernel9_Valid_Out & channel57_Kernel9_Valid_Out & channel58_Kernel9_Valid_Out & channel59_Kernel9_Valid_Out & channel60_Kernel9_Valid_Out & channel61_Kernel9_Valid_Out & channel62_Kernel9_Valid_Out & channel63_Kernel9_Valid_Out & channel64_Kernel9_Valid_Out;

	wire channel1_Kernel10_Valid_Out, channel2_Kernel10_Valid_Out, channel3_Kernel10_Valid_Out, channel4_Kernel10_Valid_Out, channel5_Kernel10_Valid_Out, channel6_Kernel10_Valid_Out, channel7_Kernel10_Valid_Out, channel8_Kernel10_Valid_Out, channel9_Kernel10_Valid_Out, channel10_Kernel10_Valid_Out, channel11_Kernel10_Valid_Out, channel12_Kernel10_Valid_Out, channel13_Kernel10_Valid_Out, channel14_Kernel10_Valid_Out, channel15_Kernel10_Valid_Out, channel16_Kernel10_Valid_Out, channel17_Kernel10_Valid_Out, channel18_Kernel10_Valid_Out, channel19_Kernel10_Valid_Out, channel20_Kernel10_Valid_Out, channel21_Kernel10_Valid_Out, channel22_Kernel10_Valid_Out, channel23_Kernel10_Valid_Out, channel24_Kernel10_Valid_Out, channel25_Kernel10_Valid_Out, channel26_Kernel10_Valid_Out, channel27_Kernel10_Valid_Out, channel28_Kernel10_Valid_Out, channel29_Kernel10_Valid_Out, channel30_Kernel10_Valid_Out, channel31_Kernel10_Valid_Out, channel32_Kernel10_Valid_Out, channel33_Kernel10_Valid_Out, channel34_Kernel10_Valid_Out, channel35_Kernel10_Valid_Out, channel36_Kernel10_Valid_Out, channel37_Kernel10_Valid_Out, channel38_Kernel10_Valid_Out, channel39_Kernel10_Valid_Out, channel40_Kernel10_Valid_Out, channel41_Kernel10_Valid_Out, channel42_Kernel10_Valid_Out, channel43_Kernel10_Valid_Out, channel44_Kernel10_Valid_Out, channel45_Kernel10_Valid_Out, channel46_Kernel10_Valid_Out, channel47_Kernel10_Valid_Out, channel48_Kernel10_Valid_Out, channel49_Kernel10_Valid_Out, channel50_Kernel10_Valid_Out, channel51_Kernel10_Valid_Out, channel52_Kernel10_Valid_Out, channel53_Kernel10_Valid_Out, channel54_Kernel10_Valid_Out, channel55_Kernel10_Valid_Out, channel56_Kernel10_Valid_Out, channel57_Kernel10_Valid_Out, channel58_Kernel10_Valid_Out, channel59_Kernel10_Valid_Out, channel60_Kernel10_Valid_Out, channel61_Kernel10_Valid_Out, channel62_Kernel10_Valid_Out, channel63_Kernel10_Valid_Out, channel64_Kernel10_Valid_Out;

	assign add_kernel10=channel1_Kernel10_Valid_Out & channel2_Kernel10_Valid_Out & channel3_Kernel10_Valid_Out & channel4_Kernel10_Valid_Out & channel5_Kernel10_Valid_Out & channel6_Kernel10_Valid_Out & channel7_Kernel10_Valid_Out & channel8_Kernel10_Valid_Out & channel9_Kernel10_Valid_Out & channel10_Kernel10_Valid_Out & channel11_Kernel10_Valid_Out & channel12_Kernel10_Valid_Out & channel13_Kernel10_Valid_Out & channel14_Kernel10_Valid_Out & channel15_Kernel10_Valid_Out & channel16_Kernel10_Valid_Out & channel17_Kernel10_Valid_Out & channel18_Kernel10_Valid_Out & channel19_Kernel10_Valid_Out & channel20_Kernel10_Valid_Out & channel21_Kernel10_Valid_Out & channel22_Kernel10_Valid_Out & channel23_Kernel10_Valid_Out & channel24_Kernel10_Valid_Out & channel25_Kernel10_Valid_Out & channel26_Kernel10_Valid_Out & channel27_Kernel10_Valid_Out & channel28_Kernel10_Valid_Out & channel29_Kernel10_Valid_Out & channel30_Kernel10_Valid_Out & channel31_Kernel10_Valid_Out & channel32_Kernel10_Valid_Out & channel33_Kernel10_Valid_Out & channel34_Kernel10_Valid_Out & channel35_Kernel10_Valid_Out & channel36_Kernel10_Valid_Out & channel37_Kernel10_Valid_Out & channel38_Kernel10_Valid_Out & channel39_Kernel10_Valid_Out & channel40_Kernel10_Valid_Out & channel41_Kernel10_Valid_Out & channel42_Kernel10_Valid_Out & channel43_Kernel10_Valid_Out & channel44_Kernel10_Valid_Out & channel45_Kernel10_Valid_Out & channel46_Kernel10_Valid_Out & channel47_Kernel10_Valid_Out & channel48_Kernel10_Valid_Out & channel49_Kernel10_Valid_Out & channel50_Kernel10_Valid_Out & channel51_Kernel10_Valid_Out & channel52_Kernel10_Valid_Out & channel53_Kernel10_Valid_Out & channel54_Kernel10_Valid_Out & channel55_Kernel10_Valid_Out & channel56_Kernel10_Valid_Out & channel57_Kernel10_Valid_Out & channel58_Kernel10_Valid_Out & channel59_Kernel10_Valid_Out & channel60_Kernel10_Valid_Out & channel61_Kernel10_Valid_Out & channel62_Kernel10_Valid_Out & channel63_Kernel10_Valid_Out & channel64_Kernel10_Valid_Out;

	wire channel1_Kernel11_Valid_Out, channel2_Kernel11_Valid_Out, channel3_Kernel11_Valid_Out, channel4_Kernel11_Valid_Out, channel5_Kernel11_Valid_Out, channel6_Kernel11_Valid_Out, channel7_Kernel11_Valid_Out, channel8_Kernel11_Valid_Out, channel9_Kernel11_Valid_Out, channel10_Kernel11_Valid_Out, channel11_Kernel11_Valid_Out, channel12_Kernel11_Valid_Out, channel13_Kernel11_Valid_Out, channel14_Kernel11_Valid_Out, channel15_Kernel11_Valid_Out, channel16_Kernel11_Valid_Out, channel17_Kernel11_Valid_Out, channel18_Kernel11_Valid_Out, channel19_Kernel11_Valid_Out, channel20_Kernel11_Valid_Out, channel21_Kernel11_Valid_Out, channel22_Kernel11_Valid_Out, channel23_Kernel11_Valid_Out, channel24_Kernel11_Valid_Out, channel25_Kernel11_Valid_Out, channel26_Kernel11_Valid_Out, channel27_Kernel11_Valid_Out, channel28_Kernel11_Valid_Out, channel29_Kernel11_Valid_Out, channel30_Kernel11_Valid_Out, channel31_Kernel11_Valid_Out, channel32_Kernel11_Valid_Out, channel33_Kernel11_Valid_Out, channel34_Kernel11_Valid_Out, channel35_Kernel11_Valid_Out, channel36_Kernel11_Valid_Out, channel37_Kernel11_Valid_Out, channel38_Kernel11_Valid_Out, channel39_Kernel11_Valid_Out, channel40_Kernel11_Valid_Out, channel41_Kernel11_Valid_Out, channel42_Kernel11_Valid_Out, channel43_Kernel11_Valid_Out, channel44_Kernel11_Valid_Out, channel45_Kernel11_Valid_Out, channel46_Kernel11_Valid_Out, channel47_Kernel11_Valid_Out, channel48_Kernel11_Valid_Out, channel49_Kernel11_Valid_Out, channel50_Kernel11_Valid_Out, channel51_Kernel11_Valid_Out, channel52_Kernel11_Valid_Out, channel53_Kernel11_Valid_Out, channel54_Kernel11_Valid_Out, channel55_Kernel11_Valid_Out, channel56_Kernel11_Valid_Out, channel57_Kernel11_Valid_Out, channel58_Kernel11_Valid_Out, channel59_Kernel11_Valid_Out, channel60_Kernel11_Valid_Out, channel61_Kernel11_Valid_Out, channel62_Kernel11_Valid_Out, channel63_Kernel11_Valid_Out, channel64_Kernel11_Valid_Out;

	assign add_kernel11=channel1_Kernel11_Valid_Out & channel2_Kernel11_Valid_Out & channel3_Kernel11_Valid_Out & channel4_Kernel11_Valid_Out & channel5_Kernel11_Valid_Out & channel6_Kernel11_Valid_Out & channel7_Kernel11_Valid_Out & channel8_Kernel11_Valid_Out & channel9_Kernel11_Valid_Out & channel10_Kernel11_Valid_Out & channel11_Kernel11_Valid_Out & channel12_Kernel11_Valid_Out & channel13_Kernel11_Valid_Out & channel14_Kernel11_Valid_Out & channel15_Kernel11_Valid_Out & channel16_Kernel11_Valid_Out & channel17_Kernel11_Valid_Out & channel18_Kernel11_Valid_Out & channel19_Kernel11_Valid_Out & channel20_Kernel11_Valid_Out & channel21_Kernel11_Valid_Out & channel22_Kernel11_Valid_Out & channel23_Kernel11_Valid_Out & channel24_Kernel11_Valid_Out & channel25_Kernel11_Valid_Out & channel26_Kernel11_Valid_Out & channel27_Kernel11_Valid_Out & channel28_Kernel11_Valid_Out & channel29_Kernel11_Valid_Out & channel30_Kernel11_Valid_Out & channel31_Kernel11_Valid_Out & channel32_Kernel11_Valid_Out & channel33_Kernel11_Valid_Out & channel34_Kernel11_Valid_Out & channel35_Kernel11_Valid_Out & channel36_Kernel11_Valid_Out & channel37_Kernel11_Valid_Out & channel38_Kernel11_Valid_Out & channel39_Kernel11_Valid_Out & channel40_Kernel11_Valid_Out & channel41_Kernel11_Valid_Out & channel42_Kernel11_Valid_Out & channel43_Kernel11_Valid_Out & channel44_Kernel11_Valid_Out & channel45_Kernel11_Valid_Out & channel46_Kernel11_Valid_Out & channel47_Kernel11_Valid_Out & channel48_Kernel11_Valid_Out & channel49_Kernel11_Valid_Out & channel50_Kernel11_Valid_Out & channel51_Kernel11_Valid_Out & channel52_Kernel11_Valid_Out & channel53_Kernel11_Valid_Out & channel54_Kernel11_Valid_Out & channel55_Kernel11_Valid_Out & channel56_Kernel11_Valid_Out & channel57_Kernel11_Valid_Out & channel58_Kernel11_Valid_Out & channel59_Kernel11_Valid_Out & channel60_Kernel11_Valid_Out & channel61_Kernel11_Valid_Out & channel62_Kernel11_Valid_Out & channel63_Kernel11_Valid_Out & channel64_Kernel11_Valid_Out;

	wire channel1_Kernel12_Valid_Out, channel2_Kernel12_Valid_Out, channel3_Kernel12_Valid_Out, channel4_Kernel12_Valid_Out, channel5_Kernel12_Valid_Out, channel6_Kernel12_Valid_Out, channel7_Kernel12_Valid_Out, channel8_Kernel12_Valid_Out, channel9_Kernel12_Valid_Out, channel10_Kernel12_Valid_Out, channel11_Kernel12_Valid_Out, channel12_Kernel12_Valid_Out, channel13_Kernel12_Valid_Out, channel14_Kernel12_Valid_Out, channel15_Kernel12_Valid_Out, channel16_Kernel12_Valid_Out, channel17_Kernel12_Valid_Out, channel18_Kernel12_Valid_Out, channel19_Kernel12_Valid_Out, channel20_Kernel12_Valid_Out, channel21_Kernel12_Valid_Out, channel22_Kernel12_Valid_Out, channel23_Kernel12_Valid_Out, channel24_Kernel12_Valid_Out, channel25_Kernel12_Valid_Out, channel26_Kernel12_Valid_Out, channel27_Kernel12_Valid_Out, channel28_Kernel12_Valid_Out, channel29_Kernel12_Valid_Out, channel30_Kernel12_Valid_Out, channel31_Kernel12_Valid_Out, channel32_Kernel12_Valid_Out, channel33_Kernel12_Valid_Out, channel34_Kernel12_Valid_Out, channel35_Kernel12_Valid_Out, channel36_Kernel12_Valid_Out, channel37_Kernel12_Valid_Out, channel38_Kernel12_Valid_Out, channel39_Kernel12_Valid_Out, channel40_Kernel12_Valid_Out, channel41_Kernel12_Valid_Out, channel42_Kernel12_Valid_Out, channel43_Kernel12_Valid_Out, channel44_Kernel12_Valid_Out, channel45_Kernel12_Valid_Out, channel46_Kernel12_Valid_Out, channel47_Kernel12_Valid_Out, channel48_Kernel12_Valid_Out, channel49_Kernel12_Valid_Out, channel50_Kernel12_Valid_Out, channel51_Kernel12_Valid_Out, channel52_Kernel12_Valid_Out, channel53_Kernel12_Valid_Out, channel54_Kernel12_Valid_Out, channel55_Kernel12_Valid_Out, channel56_Kernel12_Valid_Out, channel57_Kernel12_Valid_Out, channel58_Kernel12_Valid_Out, channel59_Kernel12_Valid_Out, channel60_Kernel12_Valid_Out, channel61_Kernel12_Valid_Out, channel62_Kernel12_Valid_Out, channel63_Kernel12_Valid_Out, channel64_Kernel12_Valid_Out;

	assign add_kernel12=channel1_Kernel12_Valid_Out & channel2_Kernel12_Valid_Out & channel3_Kernel12_Valid_Out & channel4_Kernel12_Valid_Out & channel5_Kernel12_Valid_Out & channel6_Kernel12_Valid_Out & channel7_Kernel12_Valid_Out & channel8_Kernel12_Valid_Out & channel9_Kernel12_Valid_Out & channel10_Kernel12_Valid_Out & channel11_Kernel12_Valid_Out & channel12_Kernel12_Valid_Out & channel13_Kernel12_Valid_Out & channel14_Kernel12_Valid_Out & channel15_Kernel12_Valid_Out & channel16_Kernel12_Valid_Out & channel17_Kernel12_Valid_Out & channel18_Kernel12_Valid_Out & channel19_Kernel12_Valid_Out & channel20_Kernel12_Valid_Out & channel21_Kernel12_Valid_Out & channel22_Kernel12_Valid_Out & channel23_Kernel12_Valid_Out & channel24_Kernel12_Valid_Out & channel25_Kernel12_Valid_Out & channel26_Kernel12_Valid_Out & channel27_Kernel12_Valid_Out & channel28_Kernel12_Valid_Out & channel29_Kernel12_Valid_Out & channel30_Kernel12_Valid_Out & channel31_Kernel12_Valid_Out & channel32_Kernel12_Valid_Out & channel33_Kernel12_Valid_Out & channel34_Kernel12_Valid_Out & channel35_Kernel12_Valid_Out & channel36_Kernel12_Valid_Out & channel37_Kernel12_Valid_Out & channel38_Kernel12_Valid_Out & channel39_Kernel12_Valid_Out & channel40_Kernel12_Valid_Out & channel41_Kernel12_Valid_Out & channel42_Kernel12_Valid_Out & channel43_Kernel12_Valid_Out & channel44_Kernel12_Valid_Out & channel45_Kernel12_Valid_Out & channel46_Kernel12_Valid_Out & channel47_Kernel12_Valid_Out & channel48_Kernel12_Valid_Out & channel49_Kernel12_Valid_Out & channel50_Kernel12_Valid_Out & channel51_Kernel12_Valid_Out & channel52_Kernel12_Valid_Out & channel53_Kernel12_Valid_Out & channel54_Kernel12_Valid_Out & channel55_Kernel12_Valid_Out & channel56_Kernel12_Valid_Out & channel57_Kernel12_Valid_Out & channel58_Kernel12_Valid_Out & channel59_Kernel12_Valid_Out & channel60_Kernel12_Valid_Out & channel61_Kernel12_Valid_Out & channel62_Kernel12_Valid_Out & channel63_Kernel12_Valid_Out & channel64_Kernel12_Valid_Out;

	wire channel1_Kernel13_Valid_Out, channel2_Kernel13_Valid_Out, channel3_Kernel13_Valid_Out, channel4_Kernel13_Valid_Out, channel5_Kernel13_Valid_Out, channel6_Kernel13_Valid_Out, channel7_Kernel13_Valid_Out, channel8_Kernel13_Valid_Out, channel9_Kernel13_Valid_Out, channel10_Kernel13_Valid_Out, channel11_Kernel13_Valid_Out, channel12_Kernel13_Valid_Out, channel13_Kernel13_Valid_Out, channel14_Kernel13_Valid_Out, channel15_Kernel13_Valid_Out, channel16_Kernel13_Valid_Out, channel17_Kernel13_Valid_Out, channel18_Kernel13_Valid_Out, channel19_Kernel13_Valid_Out, channel20_Kernel13_Valid_Out, channel21_Kernel13_Valid_Out, channel22_Kernel13_Valid_Out, channel23_Kernel13_Valid_Out, channel24_Kernel13_Valid_Out, channel25_Kernel13_Valid_Out, channel26_Kernel13_Valid_Out, channel27_Kernel13_Valid_Out, channel28_Kernel13_Valid_Out, channel29_Kernel13_Valid_Out, channel30_Kernel13_Valid_Out, channel31_Kernel13_Valid_Out, channel32_Kernel13_Valid_Out, channel33_Kernel13_Valid_Out, channel34_Kernel13_Valid_Out, channel35_Kernel13_Valid_Out, channel36_Kernel13_Valid_Out, channel37_Kernel13_Valid_Out, channel38_Kernel13_Valid_Out, channel39_Kernel13_Valid_Out, channel40_Kernel13_Valid_Out, channel41_Kernel13_Valid_Out, channel42_Kernel13_Valid_Out, channel43_Kernel13_Valid_Out, channel44_Kernel13_Valid_Out, channel45_Kernel13_Valid_Out, channel46_Kernel13_Valid_Out, channel47_Kernel13_Valid_Out, channel48_Kernel13_Valid_Out, channel49_Kernel13_Valid_Out, channel50_Kernel13_Valid_Out, channel51_Kernel13_Valid_Out, channel52_Kernel13_Valid_Out, channel53_Kernel13_Valid_Out, channel54_Kernel13_Valid_Out, channel55_Kernel13_Valid_Out, channel56_Kernel13_Valid_Out, channel57_Kernel13_Valid_Out, channel58_Kernel13_Valid_Out, channel59_Kernel13_Valid_Out, channel60_Kernel13_Valid_Out, channel61_Kernel13_Valid_Out, channel62_Kernel13_Valid_Out, channel63_Kernel13_Valid_Out, channel64_Kernel13_Valid_Out;

	assign add_kernel13=channel1_Kernel13_Valid_Out & channel2_Kernel13_Valid_Out & channel3_Kernel13_Valid_Out & channel4_Kernel13_Valid_Out & channel5_Kernel13_Valid_Out & channel6_Kernel13_Valid_Out & channel7_Kernel13_Valid_Out & channel8_Kernel13_Valid_Out & channel9_Kernel13_Valid_Out & channel10_Kernel13_Valid_Out & channel11_Kernel13_Valid_Out & channel12_Kernel13_Valid_Out & channel13_Kernel13_Valid_Out & channel14_Kernel13_Valid_Out & channel15_Kernel13_Valid_Out & channel16_Kernel13_Valid_Out & channel17_Kernel13_Valid_Out & channel18_Kernel13_Valid_Out & channel19_Kernel13_Valid_Out & channel20_Kernel13_Valid_Out & channel21_Kernel13_Valid_Out & channel22_Kernel13_Valid_Out & channel23_Kernel13_Valid_Out & channel24_Kernel13_Valid_Out & channel25_Kernel13_Valid_Out & channel26_Kernel13_Valid_Out & channel27_Kernel13_Valid_Out & channel28_Kernel13_Valid_Out & channel29_Kernel13_Valid_Out & channel30_Kernel13_Valid_Out & channel31_Kernel13_Valid_Out & channel32_Kernel13_Valid_Out & channel33_Kernel13_Valid_Out & channel34_Kernel13_Valid_Out & channel35_Kernel13_Valid_Out & channel36_Kernel13_Valid_Out & channel37_Kernel13_Valid_Out & channel38_Kernel13_Valid_Out & channel39_Kernel13_Valid_Out & channel40_Kernel13_Valid_Out & channel41_Kernel13_Valid_Out & channel42_Kernel13_Valid_Out & channel43_Kernel13_Valid_Out & channel44_Kernel13_Valid_Out & channel45_Kernel13_Valid_Out & channel46_Kernel13_Valid_Out & channel47_Kernel13_Valid_Out & channel48_Kernel13_Valid_Out & channel49_Kernel13_Valid_Out & channel50_Kernel13_Valid_Out & channel51_Kernel13_Valid_Out & channel52_Kernel13_Valid_Out & channel53_Kernel13_Valid_Out & channel54_Kernel13_Valid_Out & channel55_Kernel13_Valid_Out & channel56_Kernel13_Valid_Out & channel57_Kernel13_Valid_Out & channel58_Kernel13_Valid_Out & channel59_Kernel13_Valid_Out & channel60_Kernel13_Valid_Out & channel61_Kernel13_Valid_Out & channel62_Kernel13_Valid_Out & channel63_Kernel13_Valid_Out & channel64_Kernel13_Valid_Out;

	wire channel1_Kernel14_Valid_Out, channel2_Kernel14_Valid_Out, channel3_Kernel14_Valid_Out, channel4_Kernel14_Valid_Out, channel5_Kernel14_Valid_Out, channel6_Kernel14_Valid_Out, channel7_Kernel14_Valid_Out, channel8_Kernel14_Valid_Out, channel9_Kernel14_Valid_Out, channel10_Kernel14_Valid_Out, channel11_Kernel14_Valid_Out, channel12_Kernel14_Valid_Out, channel13_Kernel14_Valid_Out, channel14_Kernel14_Valid_Out, channel15_Kernel14_Valid_Out, channel16_Kernel14_Valid_Out, channel17_Kernel14_Valid_Out, channel18_Kernel14_Valid_Out, channel19_Kernel14_Valid_Out, channel20_Kernel14_Valid_Out, channel21_Kernel14_Valid_Out, channel22_Kernel14_Valid_Out, channel23_Kernel14_Valid_Out, channel24_Kernel14_Valid_Out, channel25_Kernel14_Valid_Out, channel26_Kernel14_Valid_Out, channel27_Kernel14_Valid_Out, channel28_Kernel14_Valid_Out, channel29_Kernel14_Valid_Out, channel30_Kernel14_Valid_Out, channel31_Kernel14_Valid_Out, channel32_Kernel14_Valid_Out, channel33_Kernel14_Valid_Out, channel34_Kernel14_Valid_Out, channel35_Kernel14_Valid_Out, channel36_Kernel14_Valid_Out, channel37_Kernel14_Valid_Out, channel38_Kernel14_Valid_Out, channel39_Kernel14_Valid_Out, channel40_Kernel14_Valid_Out, channel41_Kernel14_Valid_Out, channel42_Kernel14_Valid_Out, channel43_Kernel14_Valid_Out, channel44_Kernel14_Valid_Out, channel45_Kernel14_Valid_Out, channel46_Kernel14_Valid_Out, channel47_Kernel14_Valid_Out, channel48_Kernel14_Valid_Out, channel49_Kernel14_Valid_Out, channel50_Kernel14_Valid_Out, channel51_Kernel14_Valid_Out, channel52_Kernel14_Valid_Out, channel53_Kernel14_Valid_Out, channel54_Kernel14_Valid_Out, channel55_Kernel14_Valid_Out, channel56_Kernel14_Valid_Out, channel57_Kernel14_Valid_Out, channel58_Kernel14_Valid_Out, channel59_Kernel14_Valid_Out, channel60_Kernel14_Valid_Out, channel61_Kernel14_Valid_Out, channel62_Kernel14_Valid_Out, channel63_Kernel14_Valid_Out, channel64_Kernel14_Valid_Out;

	assign add_kernel14=channel1_Kernel14_Valid_Out & channel2_Kernel14_Valid_Out & channel3_Kernel14_Valid_Out & channel4_Kernel14_Valid_Out & channel5_Kernel14_Valid_Out & channel6_Kernel14_Valid_Out & channel7_Kernel14_Valid_Out & channel8_Kernel14_Valid_Out & channel9_Kernel14_Valid_Out & channel10_Kernel14_Valid_Out & channel11_Kernel14_Valid_Out & channel12_Kernel14_Valid_Out & channel13_Kernel14_Valid_Out & channel14_Kernel14_Valid_Out & channel15_Kernel14_Valid_Out & channel16_Kernel14_Valid_Out & channel17_Kernel14_Valid_Out & channel18_Kernel14_Valid_Out & channel19_Kernel14_Valid_Out & channel20_Kernel14_Valid_Out & channel21_Kernel14_Valid_Out & channel22_Kernel14_Valid_Out & channel23_Kernel14_Valid_Out & channel24_Kernel14_Valid_Out & channel25_Kernel14_Valid_Out & channel26_Kernel14_Valid_Out & channel27_Kernel14_Valid_Out & channel28_Kernel14_Valid_Out & channel29_Kernel14_Valid_Out & channel30_Kernel14_Valid_Out & channel31_Kernel14_Valid_Out & channel32_Kernel14_Valid_Out & channel33_Kernel14_Valid_Out & channel34_Kernel14_Valid_Out & channel35_Kernel14_Valid_Out & channel36_Kernel14_Valid_Out & channel37_Kernel14_Valid_Out & channel38_Kernel14_Valid_Out & channel39_Kernel14_Valid_Out & channel40_Kernel14_Valid_Out & channel41_Kernel14_Valid_Out & channel42_Kernel14_Valid_Out & channel43_Kernel14_Valid_Out & channel44_Kernel14_Valid_Out & channel45_Kernel14_Valid_Out & channel46_Kernel14_Valid_Out & channel47_Kernel14_Valid_Out & channel48_Kernel14_Valid_Out & channel49_Kernel14_Valid_Out & channel50_Kernel14_Valid_Out & channel51_Kernel14_Valid_Out & channel52_Kernel14_Valid_Out & channel53_Kernel14_Valid_Out & channel54_Kernel14_Valid_Out & channel55_Kernel14_Valid_Out & channel56_Kernel14_Valid_Out & channel57_Kernel14_Valid_Out & channel58_Kernel14_Valid_Out & channel59_Kernel14_Valid_Out & channel60_Kernel14_Valid_Out & channel61_Kernel14_Valid_Out & channel62_Kernel14_Valid_Out & channel63_Kernel14_Valid_Out & channel64_Kernel14_Valid_Out;

	wire channel1_Kernel15_Valid_Out, channel2_Kernel15_Valid_Out, channel3_Kernel15_Valid_Out, channel4_Kernel15_Valid_Out, channel5_Kernel15_Valid_Out, channel6_Kernel15_Valid_Out, channel7_Kernel15_Valid_Out, channel8_Kernel15_Valid_Out, channel9_Kernel15_Valid_Out, channel10_Kernel15_Valid_Out, channel11_Kernel15_Valid_Out, channel12_Kernel15_Valid_Out, channel13_Kernel15_Valid_Out, channel14_Kernel15_Valid_Out, channel15_Kernel15_Valid_Out, channel16_Kernel15_Valid_Out, channel17_Kernel15_Valid_Out, channel18_Kernel15_Valid_Out, channel19_Kernel15_Valid_Out, channel20_Kernel15_Valid_Out, channel21_Kernel15_Valid_Out, channel22_Kernel15_Valid_Out, channel23_Kernel15_Valid_Out, channel24_Kernel15_Valid_Out, channel25_Kernel15_Valid_Out, channel26_Kernel15_Valid_Out, channel27_Kernel15_Valid_Out, channel28_Kernel15_Valid_Out, channel29_Kernel15_Valid_Out, channel30_Kernel15_Valid_Out, channel31_Kernel15_Valid_Out, channel32_Kernel15_Valid_Out, channel33_Kernel15_Valid_Out, channel34_Kernel15_Valid_Out, channel35_Kernel15_Valid_Out, channel36_Kernel15_Valid_Out, channel37_Kernel15_Valid_Out, channel38_Kernel15_Valid_Out, channel39_Kernel15_Valid_Out, channel40_Kernel15_Valid_Out, channel41_Kernel15_Valid_Out, channel42_Kernel15_Valid_Out, channel43_Kernel15_Valid_Out, channel44_Kernel15_Valid_Out, channel45_Kernel15_Valid_Out, channel46_Kernel15_Valid_Out, channel47_Kernel15_Valid_Out, channel48_Kernel15_Valid_Out, channel49_Kernel15_Valid_Out, channel50_Kernel15_Valid_Out, channel51_Kernel15_Valid_Out, channel52_Kernel15_Valid_Out, channel53_Kernel15_Valid_Out, channel54_Kernel15_Valid_Out, channel55_Kernel15_Valid_Out, channel56_Kernel15_Valid_Out, channel57_Kernel15_Valid_Out, channel58_Kernel15_Valid_Out, channel59_Kernel15_Valid_Out, channel60_Kernel15_Valid_Out, channel61_Kernel15_Valid_Out, channel62_Kernel15_Valid_Out, channel63_Kernel15_Valid_Out, channel64_Kernel15_Valid_Out;

	assign add_kernel15=channel1_Kernel15_Valid_Out & channel2_Kernel15_Valid_Out & channel3_Kernel15_Valid_Out & channel4_Kernel15_Valid_Out & channel5_Kernel15_Valid_Out & channel6_Kernel15_Valid_Out & channel7_Kernel15_Valid_Out & channel8_Kernel15_Valid_Out & channel9_Kernel15_Valid_Out & channel10_Kernel15_Valid_Out & channel11_Kernel15_Valid_Out & channel12_Kernel15_Valid_Out & channel13_Kernel15_Valid_Out & channel14_Kernel15_Valid_Out & channel15_Kernel15_Valid_Out & channel16_Kernel15_Valid_Out & channel17_Kernel15_Valid_Out & channel18_Kernel15_Valid_Out & channel19_Kernel15_Valid_Out & channel20_Kernel15_Valid_Out & channel21_Kernel15_Valid_Out & channel22_Kernel15_Valid_Out & channel23_Kernel15_Valid_Out & channel24_Kernel15_Valid_Out & channel25_Kernel15_Valid_Out & channel26_Kernel15_Valid_Out & channel27_Kernel15_Valid_Out & channel28_Kernel15_Valid_Out & channel29_Kernel15_Valid_Out & channel30_Kernel15_Valid_Out & channel31_Kernel15_Valid_Out & channel32_Kernel15_Valid_Out & channel33_Kernel15_Valid_Out & channel34_Kernel15_Valid_Out & channel35_Kernel15_Valid_Out & channel36_Kernel15_Valid_Out & channel37_Kernel15_Valid_Out & channel38_Kernel15_Valid_Out & channel39_Kernel15_Valid_Out & channel40_Kernel15_Valid_Out & channel41_Kernel15_Valid_Out & channel42_Kernel15_Valid_Out & channel43_Kernel15_Valid_Out & channel44_Kernel15_Valid_Out & channel45_Kernel15_Valid_Out & channel46_Kernel15_Valid_Out & channel47_Kernel15_Valid_Out & channel48_Kernel15_Valid_Out & channel49_Kernel15_Valid_Out & channel50_Kernel15_Valid_Out & channel51_Kernel15_Valid_Out & channel52_Kernel15_Valid_Out & channel53_Kernel15_Valid_Out & channel54_Kernel15_Valid_Out & channel55_Kernel15_Valid_Out & channel56_Kernel15_Valid_Out & channel57_Kernel15_Valid_Out & channel58_Kernel15_Valid_Out & channel59_Kernel15_Valid_Out & channel60_Kernel15_Valid_Out & channel61_Kernel15_Valid_Out & channel62_Kernel15_Valid_Out & channel63_Kernel15_Valid_Out & channel64_Kernel15_Valid_Out;

	wire channel1_Kernel16_Valid_Out, channel2_Kernel16_Valid_Out, channel3_Kernel16_Valid_Out, channel4_Kernel16_Valid_Out, channel5_Kernel16_Valid_Out, channel6_Kernel16_Valid_Out, channel7_Kernel16_Valid_Out, channel8_Kernel16_Valid_Out, channel9_Kernel16_Valid_Out, channel10_Kernel16_Valid_Out, channel11_Kernel16_Valid_Out, channel12_Kernel16_Valid_Out, channel13_Kernel16_Valid_Out, channel14_Kernel16_Valid_Out, channel15_Kernel16_Valid_Out, channel16_Kernel16_Valid_Out, channel17_Kernel16_Valid_Out, channel18_Kernel16_Valid_Out, channel19_Kernel16_Valid_Out, channel20_Kernel16_Valid_Out, channel21_Kernel16_Valid_Out, channel22_Kernel16_Valid_Out, channel23_Kernel16_Valid_Out, channel24_Kernel16_Valid_Out, channel25_Kernel16_Valid_Out, channel26_Kernel16_Valid_Out, channel27_Kernel16_Valid_Out, channel28_Kernel16_Valid_Out, channel29_Kernel16_Valid_Out, channel30_Kernel16_Valid_Out, channel31_Kernel16_Valid_Out, channel32_Kernel16_Valid_Out, channel33_Kernel16_Valid_Out, channel34_Kernel16_Valid_Out, channel35_Kernel16_Valid_Out, channel36_Kernel16_Valid_Out, channel37_Kernel16_Valid_Out, channel38_Kernel16_Valid_Out, channel39_Kernel16_Valid_Out, channel40_Kernel16_Valid_Out, channel41_Kernel16_Valid_Out, channel42_Kernel16_Valid_Out, channel43_Kernel16_Valid_Out, channel44_Kernel16_Valid_Out, channel45_Kernel16_Valid_Out, channel46_Kernel16_Valid_Out, channel47_Kernel16_Valid_Out, channel48_Kernel16_Valid_Out, channel49_Kernel16_Valid_Out, channel50_Kernel16_Valid_Out, channel51_Kernel16_Valid_Out, channel52_Kernel16_Valid_Out, channel53_Kernel16_Valid_Out, channel54_Kernel16_Valid_Out, channel55_Kernel16_Valid_Out, channel56_Kernel16_Valid_Out, channel57_Kernel16_Valid_Out, channel58_Kernel16_Valid_Out, channel59_Kernel16_Valid_Out, channel60_Kernel16_Valid_Out, channel61_Kernel16_Valid_Out, channel62_Kernel16_Valid_Out, channel63_Kernel16_Valid_Out, channel64_Kernel16_Valid_Out;

	assign add_kernel16=channel1_Kernel16_Valid_Out & channel2_Kernel16_Valid_Out & channel3_Kernel16_Valid_Out & channel4_Kernel16_Valid_Out & channel5_Kernel16_Valid_Out & channel6_Kernel16_Valid_Out & channel7_Kernel16_Valid_Out & channel8_Kernel16_Valid_Out & channel9_Kernel16_Valid_Out & channel10_Kernel16_Valid_Out & channel11_Kernel16_Valid_Out & channel12_Kernel16_Valid_Out & channel13_Kernel16_Valid_Out & channel14_Kernel16_Valid_Out & channel15_Kernel16_Valid_Out & channel16_Kernel16_Valid_Out & channel17_Kernel16_Valid_Out & channel18_Kernel16_Valid_Out & channel19_Kernel16_Valid_Out & channel20_Kernel16_Valid_Out & channel21_Kernel16_Valid_Out & channel22_Kernel16_Valid_Out & channel23_Kernel16_Valid_Out & channel24_Kernel16_Valid_Out & channel25_Kernel16_Valid_Out & channel26_Kernel16_Valid_Out & channel27_Kernel16_Valid_Out & channel28_Kernel16_Valid_Out & channel29_Kernel16_Valid_Out & channel30_Kernel16_Valid_Out & channel31_Kernel16_Valid_Out & channel32_Kernel16_Valid_Out & channel33_Kernel16_Valid_Out & channel34_Kernel16_Valid_Out & channel35_Kernel16_Valid_Out & channel36_Kernel16_Valid_Out & channel37_Kernel16_Valid_Out & channel38_Kernel16_Valid_Out & channel39_Kernel16_Valid_Out & channel40_Kernel16_Valid_Out & channel41_Kernel16_Valid_Out & channel42_Kernel16_Valid_Out & channel43_Kernel16_Valid_Out & channel44_Kernel16_Valid_Out & channel45_Kernel16_Valid_Out & channel46_Kernel16_Valid_Out & channel47_Kernel16_Valid_Out & channel48_Kernel16_Valid_Out & channel49_Kernel16_Valid_Out & channel50_Kernel16_Valid_Out & channel51_Kernel16_Valid_Out & channel52_Kernel16_Valid_Out & channel53_Kernel16_Valid_Out & channel54_Kernel16_Valid_Out & channel55_Kernel16_Valid_Out & channel56_Kernel16_Valid_Out & channel57_Kernel16_Valid_Out & channel58_Kernel16_Valid_Out & channel59_Kernel16_Valid_Out & channel60_Kernel16_Valid_Out & channel61_Kernel16_Valid_Out & channel62_Kernel16_Valid_Out & channel63_Kernel16_Valid_Out & channel64_Kernel16_Valid_Out;

	wire channel1_Kernel17_Valid_Out, channel2_Kernel17_Valid_Out, channel3_Kernel17_Valid_Out, channel4_Kernel17_Valid_Out, channel5_Kernel17_Valid_Out, channel6_Kernel17_Valid_Out, channel7_Kernel17_Valid_Out, channel8_Kernel17_Valid_Out, channel9_Kernel17_Valid_Out, channel10_Kernel17_Valid_Out, channel11_Kernel17_Valid_Out, channel12_Kernel17_Valid_Out, channel13_Kernel17_Valid_Out, channel14_Kernel17_Valid_Out, channel15_Kernel17_Valid_Out, channel16_Kernel17_Valid_Out, channel17_Kernel17_Valid_Out, channel18_Kernel17_Valid_Out, channel19_Kernel17_Valid_Out, channel20_Kernel17_Valid_Out, channel21_Kernel17_Valid_Out, channel22_Kernel17_Valid_Out, channel23_Kernel17_Valid_Out, channel24_Kernel17_Valid_Out, channel25_Kernel17_Valid_Out, channel26_Kernel17_Valid_Out, channel27_Kernel17_Valid_Out, channel28_Kernel17_Valid_Out, channel29_Kernel17_Valid_Out, channel30_Kernel17_Valid_Out, channel31_Kernel17_Valid_Out, channel32_Kernel17_Valid_Out, channel33_Kernel17_Valid_Out, channel34_Kernel17_Valid_Out, channel35_Kernel17_Valid_Out, channel36_Kernel17_Valid_Out, channel37_Kernel17_Valid_Out, channel38_Kernel17_Valid_Out, channel39_Kernel17_Valid_Out, channel40_Kernel17_Valid_Out, channel41_Kernel17_Valid_Out, channel42_Kernel17_Valid_Out, channel43_Kernel17_Valid_Out, channel44_Kernel17_Valid_Out, channel45_Kernel17_Valid_Out, channel46_Kernel17_Valid_Out, channel47_Kernel17_Valid_Out, channel48_Kernel17_Valid_Out, channel49_Kernel17_Valid_Out, channel50_Kernel17_Valid_Out, channel51_Kernel17_Valid_Out, channel52_Kernel17_Valid_Out, channel53_Kernel17_Valid_Out, channel54_Kernel17_Valid_Out, channel55_Kernel17_Valid_Out, channel56_Kernel17_Valid_Out, channel57_Kernel17_Valid_Out, channel58_Kernel17_Valid_Out, channel59_Kernel17_Valid_Out, channel60_Kernel17_Valid_Out, channel61_Kernel17_Valid_Out, channel62_Kernel17_Valid_Out, channel63_Kernel17_Valid_Out, channel64_Kernel17_Valid_Out;

	assign add_kernel17=channel1_Kernel17_Valid_Out & channel2_Kernel17_Valid_Out & channel3_Kernel17_Valid_Out & channel4_Kernel17_Valid_Out & channel5_Kernel17_Valid_Out & channel6_Kernel17_Valid_Out & channel7_Kernel17_Valid_Out & channel8_Kernel17_Valid_Out & channel9_Kernel17_Valid_Out & channel10_Kernel17_Valid_Out & channel11_Kernel17_Valid_Out & channel12_Kernel17_Valid_Out & channel13_Kernel17_Valid_Out & channel14_Kernel17_Valid_Out & channel15_Kernel17_Valid_Out & channel16_Kernel17_Valid_Out & channel17_Kernel17_Valid_Out & channel18_Kernel17_Valid_Out & channel19_Kernel17_Valid_Out & channel20_Kernel17_Valid_Out & channel21_Kernel17_Valid_Out & channel22_Kernel17_Valid_Out & channel23_Kernel17_Valid_Out & channel24_Kernel17_Valid_Out & channel25_Kernel17_Valid_Out & channel26_Kernel17_Valid_Out & channel27_Kernel17_Valid_Out & channel28_Kernel17_Valid_Out & channel29_Kernel17_Valid_Out & channel30_Kernel17_Valid_Out & channel31_Kernel17_Valid_Out & channel32_Kernel17_Valid_Out & channel33_Kernel17_Valid_Out & channel34_Kernel17_Valid_Out & channel35_Kernel17_Valid_Out & channel36_Kernel17_Valid_Out & channel37_Kernel17_Valid_Out & channel38_Kernel17_Valid_Out & channel39_Kernel17_Valid_Out & channel40_Kernel17_Valid_Out & channel41_Kernel17_Valid_Out & channel42_Kernel17_Valid_Out & channel43_Kernel17_Valid_Out & channel44_Kernel17_Valid_Out & channel45_Kernel17_Valid_Out & channel46_Kernel17_Valid_Out & channel47_Kernel17_Valid_Out & channel48_Kernel17_Valid_Out & channel49_Kernel17_Valid_Out & channel50_Kernel17_Valid_Out & channel51_Kernel17_Valid_Out & channel52_Kernel17_Valid_Out & channel53_Kernel17_Valid_Out & channel54_Kernel17_Valid_Out & channel55_Kernel17_Valid_Out & channel56_Kernel17_Valid_Out & channel57_Kernel17_Valid_Out & channel58_Kernel17_Valid_Out & channel59_Kernel17_Valid_Out & channel60_Kernel17_Valid_Out & channel61_Kernel17_Valid_Out & channel62_Kernel17_Valid_Out & channel63_Kernel17_Valid_Out & channel64_Kernel17_Valid_Out;

	wire channel1_Kernel18_Valid_Out, channel2_Kernel18_Valid_Out, channel3_Kernel18_Valid_Out, channel4_Kernel18_Valid_Out, channel5_Kernel18_Valid_Out, channel6_Kernel18_Valid_Out, channel7_Kernel18_Valid_Out, channel8_Kernel18_Valid_Out, channel9_Kernel18_Valid_Out, channel10_Kernel18_Valid_Out, channel11_Kernel18_Valid_Out, channel12_Kernel18_Valid_Out, channel13_Kernel18_Valid_Out, channel14_Kernel18_Valid_Out, channel15_Kernel18_Valid_Out, channel16_Kernel18_Valid_Out, channel17_Kernel18_Valid_Out, channel18_Kernel18_Valid_Out, channel19_Kernel18_Valid_Out, channel20_Kernel18_Valid_Out, channel21_Kernel18_Valid_Out, channel22_Kernel18_Valid_Out, channel23_Kernel18_Valid_Out, channel24_Kernel18_Valid_Out, channel25_Kernel18_Valid_Out, channel26_Kernel18_Valid_Out, channel27_Kernel18_Valid_Out, channel28_Kernel18_Valid_Out, channel29_Kernel18_Valid_Out, channel30_Kernel18_Valid_Out, channel31_Kernel18_Valid_Out, channel32_Kernel18_Valid_Out, channel33_Kernel18_Valid_Out, channel34_Kernel18_Valid_Out, channel35_Kernel18_Valid_Out, channel36_Kernel18_Valid_Out, channel37_Kernel18_Valid_Out, channel38_Kernel18_Valid_Out, channel39_Kernel18_Valid_Out, channel40_Kernel18_Valid_Out, channel41_Kernel18_Valid_Out, channel42_Kernel18_Valid_Out, channel43_Kernel18_Valid_Out, channel44_Kernel18_Valid_Out, channel45_Kernel18_Valid_Out, channel46_Kernel18_Valid_Out, channel47_Kernel18_Valid_Out, channel48_Kernel18_Valid_Out, channel49_Kernel18_Valid_Out, channel50_Kernel18_Valid_Out, channel51_Kernel18_Valid_Out, channel52_Kernel18_Valid_Out, channel53_Kernel18_Valid_Out, channel54_Kernel18_Valid_Out, channel55_Kernel18_Valid_Out, channel56_Kernel18_Valid_Out, channel57_Kernel18_Valid_Out, channel58_Kernel18_Valid_Out, channel59_Kernel18_Valid_Out, channel60_Kernel18_Valid_Out, channel61_Kernel18_Valid_Out, channel62_Kernel18_Valid_Out, channel63_Kernel18_Valid_Out, channel64_Kernel18_Valid_Out;

	assign add_kernel18=channel1_Kernel18_Valid_Out & channel2_Kernel18_Valid_Out & channel3_Kernel18_Valid_Out & channel4_Kernel18_Valid_Out & channel5_Kernel18_Valid_Out & channel6_Kernel18_Valid_Out & channel7_Kernel18_Valid_Out & channel8_Kernel18_Valid_Out & channel9_Kernel18_Valid_Out & channel10_Kernel18_Valid_Out & channel11_Kernel18_Valid_Out & channel12_Kernel18_Valid_Out & channel13_Kernel18_Valid_Out & channel14_Kernel18_Valid_Out & channel15_Kernel18_Valid_Out & channel16_Kernel18_Valid_Out & channel17_Kernel18_Valid_Out & channel18_Kernel18_Valid_Out & channel19_Kernel18_Valid_Out & channel20_Kernel18_Valid_Out & channel21_Kernel18_Valid_Out & channel22_Kernel18_Valid_Out & channel23_Kernel18_Valid_Out & channel24_Kernel18_Valid_Out & channel25_Kernel18_Valid_Out & channel26_Kernel18_Valid_Out & channel27_Kernel18_Valid_Out & channel28_Kernel18_Valid_Out & channel29_Kernel18_Valid_Out & channel30_Kernel18_Valid_Out & channel31_Kernel18_Valid_Out & channel32_Kernel18_Valid_Out & channel33_Kernel18_Valid_Out & channel34_Kernel18_Valid_Out & channel35_Kernel18_Valid_Out & channel36_Kernel18_Valid_Out & channel37_Kernel18_Valid_Out & channel38_Kernel18_Valid_Out & channel39_Kernel18_Valid_Out & channel40_Kernel18_Valid_Out & channel41_Kernel18_Valid_Out & channel42_Kernel18_Valid_Out & channel43_Kernel18_Valid_Out & channel44_Kernel18_Valid_Out & channel45_Kernel18_Valid_Out & channel46_Kernel18_Valid_Out & channel47_Kernel18_Valid_Out & channel48_Kernel18_Valid_Out & channel49_Kernel18_Valid_Out & channel50_Kernel18_Valid_Out & channel51_Kernel18_Valid_Out & channel52_Kernel18_Valid_Out & channel53_Kernel18_Valid_Out & channel54_Kernel18_Valid_Out & channel55_Kernel18_Valid_Out & channel56_Kernel18_Valid_Out & channel57_Kernel18_Valid_Out & channel58_Kernel18_Valid_Out & channel59_Kernel18_Valid_Out & channel60_Kernel18_Valid_Out & channel61_Kernel18_Valid_Out & channel62_Kernel18_Valid_Out & channel63_Kernel18_Valid_Out & channel64_Kernel18_Valid_Out;

	wire channel1_Kernel19_Valid_Out, channel2_Kernel19_Valid_Out, channel3_Kernel19_Valid_Out, channel4_Kernel19_Valid_Out, channel5_Kernel19_Valid_Out, channel6_Kernel19_Valid_Out, channel7_Kernel19_Valid_Out, channel8_Kernel19_Valid_Out, channel9_Kernel19_Valid_Out, channel10_Kernel19_Valid_Out, channel11_Kernel19_Valid_Out, channel12_Kernel19_Valid_Out, channel13_Kernel19_Valid_Out, channel14_Kernel19_Valid_Out, channel15_Kernel19_Valid_Out, channel16_Kernel19_Valid_Out, channel17_Kernel19_Valid_Out, channel18_Kernel19_Valid_Out, channel19_Kernel19_Valid_Out, channel20_Kernel19_Valid_Out, channel21_Kernel19_Valid_Out, channel22_Kernel19_Valid_Out, channel23_Kernel19_Valid_Out, channel24_Kernel19_Valid_Out, channel25_Kernel19_Valid_Out, channel26_Kernel19_Valid_Out, channel27_Kernel19_Valid_Out, channel28_Kernel19_Valid_Out, channel29_Kernel19_Valid_Out, channel30_Kernel19_Valid_Out, channel31_Kernel19_Valid_Out, channel32_Kernel19_Valid_Out, channel33_Kernel19_Valid_Out, channel34_Kernel19_Valid_Out, channel35_Kernel19_Valid_Out, channel36_Kernel19_Valid_Out, channel37_Kernel19_Valid_Out, channel38_Kernel19_Valid_Out, channel39_Kernel19_Valid_Out, channel40_Kernel19_Valid_Out, channel41_Kernel19_Valid_Out, channel42_Kernel19_Valid_Out, channel43_Kernel19_Valid_Out, channel44_Kernel19_Valid_Out, channel45_Kernel19_Valid_Out, channel46_Kernel19_Valid_Out, channel47_Kernel19_Valid_Out, channel48_Kernel19_Valid_Out, channel49_Kernel19_Valid_Out, channel50_Kernel19_Valid_Out, channel51_Kernel19_Valid_Out, channel52_Kernel19_Valid_Out, channel53_Kernel19_Valid_Out, channel54_Kernel19_Valid_Out, channel55_Kernel19_Valid_Out, channel56_Kernel19_Valid_Out, channel57_Kernel19_Valid_Out, channel58_Kernel19_Valid_Out, channel59_Kernel19_Valid_Out, channel60_Kernel19_Valid_Out, channel61_Kernel19_Valid_Out, channel62_Kernel19_Valid_Out, channel63_Kernel19_Valid_Out, channel64_Kernel19_Valid_Out;

	assign add_kernel19=channel1_Kernel19_Valid_Out & channel2_Kernel19_Valid_Out & channel3_Kernel19_Valid_Out & channel4_Kernel19_Valid_Out & channel5_Kernel19_Valid_Out & channel6_Kernel19_Valid_Out & channel7_Kernel19_Valid_Out & channel8_Kernel19_Valid_Out & channel9_Kernel19_Valid_Out & channel10_Kernel19_Valid_Out & channel11_Kernel19_Valid_Out & channel12_Kernel19_Valid_Out & channel13_Kernel19_Valid_Out & channel14_Kernel19_Valid_Out & channel15_Kernel19_Valid_Out & channel16_Kernel19_Valid_Out & channel17_Kernel19_Valid_Out & channel18_Kernel19_Valid_Out & channel19_Kernel19_Valid_Out & channel20_Kernel19_Valid_Out & channel21_Kernel19_Valid_Out & channel22_Kernel19_Valid_Out & channel23_Kernel19_Valid_Out & channel24_Kernel19_Valid_Out & channel25_Kernel19_Valid_Out & channel26_Kernel19_Valid_Out & channel27_Kernel19_Valid_Out & channel28_Kernel19_Valid_Out & channel29_Kernel19_Valid_Out & channel30_Kernel19_Valid_Out & channel31_Kernel19_Valid_Out & channel32_Kernel19_Valid_Out & channel33_Kernel19_Valid_Out & channel34_Kernel19_Valid_Out & channel35_Kernel19_Valid_Out & channel36_Kernel19_Valid_Out & channel37_Kernel19_Valid_Out & channel38_Kernel19_Valid_Out & channel39_Kernel19_Valid_Out & channel40_Kernel19_Valid_Out & channel41_Kernel19_Valid_Out & channel42_Kernel19_Valid_Out & channel43_Kernel19_Valid_Out & channel44_Kernel19_Valid_Out & channel45_Kernel19_Valid_Out & channel46_Kernel19_Valid_Out & channel47_Kernel19_Valid_Out & channel48_Kernel19_Valid_Out & channel49_Kernel19_Valid_Out & channel50_Kernel19_Valid_Out & channel51_Kernel19_Valid_Out & channel52_Kernel19_Valid_Out & channel53_Kernel19_Valid_Out & channel54_Kernel19_Valid_Out & channel55_Kernel19_Valid_Out & channel56_Kernel19_Valid_Out & channel57_Kernel19_Valid_Out & channel58_Kernel19_Valid_Out & channel59_Kernel19_Valid_Out & channel60_Kernel19_Valid_Out & channel61_Kernel19_Valid_Out & channel62_Kernel19_Valid_Out & channel63_Kernel19_Valid_Out & channel64_Kernel19_Valid_Out;

	wire channel1_Kernel20_Valid_Out, channel2_Kernel20_Valid_Out, channel3_Kernel20_Valid_Out, channel4_Kernel20_Valid_Out, channel5_Kernel20_Valid_Out, channel6_Kernel20_Valid_Out, channel7_Kernel20_Valid_Out, channel8_Kernel20_Valid_Out, channel9_Kernel20_Valid_Out, channel10_Kernel20_Valid_Out, channel11_Kernel20_Valid_Out, channel12_Kernel20_Valid_Out, channel13_Kernel20_Valid_Out, channel14_Kernel20_Valid_Out, channel15_Kernel20_Valid_Out, channel16_Kernel20_Valid_Out, channel17_Kernel20_Valid_Out, channel18_Kernel20_Valid_Out, channel19_Kernel20_Valid_Out, channel20_Kernel20_Valid_Out, channel21_Kernel20_Valid_Out, channel22_Kernel20_Valid_Out, channel23_Kernel20_Valid_Out, channel24_Kernel20_Valid_Out, channel25_Kernel20_Valid_Out, channel26_Kernel20_Valid_Out, channel27_Kernel20_Valid_Out, channel28_Kernel20_Valid_Out, channel29_Kernel20_Valid_Out, channel30_Kernel20_Valid_Out, channel31_Kernel20_Valid_Out, channel32_Kernel20_Valid_Out, channel33_Kernel20_Valid_Out, channel34_Kernel20_Valid_Out, channel35_Kernel20_Valid_Out, channel36_Kernel20_Valid_Out, channel37_Kernel20_Valid_Out, channel38_Kernel20_Valid_Out, channel39_Kernel20_Valid_Out, channel40_Kernel20_Valid_Out, channel41_Kernel20_Valid_Out, channel42_Kernel20_Valid_Out, channel43_Kernel20_Valid_Out, channel44_Kernel20_Valid_Out, channel45_Kernel20_Valid_Out, channel46_Kernel20_Valid_Out, channel47_Kernel20_Valid_Out, channel48_Kernel20_Valid_Out, channel49_Kernel20_Valid_Out, channel50_Kernel20_Valid_Out, channel51_Kernel20_Valid_Out, channel52_Kernel20_Valid_Out, channel53_Kernel20_Valid_Out, channel54_Kernel20_Valid_Out, channel55_Kernel20_Valid_Out, channel56_Kernel20_Valid_Out, channel57_Kernel20_Valid_Out, channel58_Kernel20_Valid_Out, channel59_Kernel20_Valid_Out, channel60_Kernel20_Valid_Out, channel61_Kernel20_Valid_Out, channel62_Kernel20_Valid_Out, channel63_Kernel20_Valid_Out, channel64_Kernel20_Valid_Out;

	assign add_kernel20=channel1_Kernel20_Valid_Out & channel2_Kernel20_Valid_Out & channel3_Kernel20_Valid_Out & channel4_Kernel20_Valid_Out & channel5_Kernel20_Valid_Out & channel6_Kernel20_Valid_Out & channel7_Kernel20_Valid_Out & channel8_Kernel20_Valid_Out & channel9_Kernel20_Valid_Out & channel10_Kernel20_Valid_Out & channel11_Kernel20_Valid_Out & channel12_Kernel20_Valid_Out & channel13_Kernel20_Valid_Out & channel14_Kernel20_Valid_Out & channel15_Kernel20_Valid_Out & channel16_Kernel20_Valid_Out & channel17_Kernel20_Valid_Out & channel18_Kernel20_Valid_Out & channel19_Kernel20_Valid_Out & channel20_Kernel20_Valid_Out & channel21_Kernel20_Valid_Out & channel22_Kernel20_Valid_Out & channel23_Kernel20_Valid_Out & channel24_Kernel20_Valid_Out & channel25_Kernel20_Valid_Out & channel26_Kernel20_Valid_Out & channel27_Kernel20_Valid_Out & channel28_Kernel20_Valid_Out & channel29_Kernel20_Valid_Out & channel30_Kernel20_Valid_Out & channel31_Kernel20_Valid_Out & channel32_Kernel20_Valid_Out & channel33_Kernel20_Valid_Out & channel34_Kernel20_Valid_Out & channel35_Kernel20_Valid_Out & channel36_Kernel20_Valid_Out & channel37_Kernel20_Valid_Out & channel38_Kernel20_Valid_Out & channel39_Kernel20_Valid_Out & channel40_Kernel20_Valid_Out & channel41_Kernel20_Valid_Out & channel42_Kernel20_Valid_Out & channel43_Kernel20_Valid_Out & channel44_Kernel20_Valid_Out & channel45_Kernel20_Valid_Out & channel46_Kernel20_Valid_Out & channel47_Kernel20_Valid_Out & channel48_Kernel20_Valid_Out & channel49_Kernel20_Valid_Out & channel50_Kernel20_Valid_Out & channel51_Kernel20_Valid_Out & channel52_Kernel20_Valid_Out & channel53_Kernel20_Valid_Out & channel54_Kernel20_Valid_Out & channel55_Kernel20_Valid_Out & channel56_Kernel20_Valid_Out & channel57_Kernel20_Valid_Out & channel58_Kernel20_Valid_Out & channel59_Kernel20_Valid_Out & channel60_Kernel20_Valid_Out & channel61_Kernel20_Valid_Out & channel62_Kernel20_Valid_Out & channel63_Kernel20_Valid_Out & channel64_Kernel20_Valid_Out;

	wire channel1_Kernel21_Valid_Out, channel2_Kernel21_Valid_Out, channel3_Kernel21_Valid_Out, channel4_Kernel21_Valid_Out, channel5_Kernel21_Valid_Out, channel6_Kernel21_Valid_Out, channel7_Kernel21_Valid_Out, channel8_Kernel21_Valid_Out, channel9_Kernel21_Valid_Out, channel10_Kernel21_Valid_Out, channel11_Kernel21_Valid_Out, channel12_Kernel21_Valid_Out, channel13_Kernel21_Valid_Out, channel14_Kernel21_Valid_Out, channel15_Kernel21_Valid_Out, channel16_Kernel21_Valid_Out, channel17_Kernel21_Valid_Out, channel18_Kernel21_Valid_Out, channel19_Kernel21_Valid_Out, channel20_Kernel21_Valid_Out, channel21_Kernel21_Valid_Out, channel22_Kernel21_Valid_Out, channel23_Kernel21_Valid_Out, channel24_Kernel21_Valid_Out, channel25_Kernel21_Valid_Out, channel26_Kernel21_Valid_Out, channel27_Kernel21_Valid_Out, channel28_Kernel21_Valid_Out, channel29_Kernel21_Valid_Out, channel30_Kernel21_Valid_Out, channel31_Kernel21_Valid_Out, channel32_Kernel21_Valid_Out, channel33_Kernel21_Valid_Out, channel34_Kernel21_Valid_Out, channel35_Kernel21_Valid_Out, channel36_Kernel21_Valid_Out, channel37_Kernel21_Valid_Out, channel38_Kernel21_Valid_Out, channel39_Kernel21_Valid_Out, channel40_Kernel21_Valid_Out, channel41_Kernel21_Valid_Out, channel42_Kernel21_Valid_Out, channel43_Kernel21_Valid_Out, channel44_Kernel21_Valid_Out, channel45_Kernel21_Valid_Out, channel46_Kernel21_Valid_Out, channel47_Kernel21_Valid_Out, channel48_Kernel21_Valid_Out, channel49_Kernel21_Valid_Out, channel50_Kernel21_Valid_Out, channel51_Kernel21_Valid_Out, channel52_Kernel21_Valid_Out, channel53_Kernel21_Valid_Out, channel54_Kernel21_Valid_Out, channel55_Kernel21_Valid_Out, channel56_Kernel21_Valid_Out, channel57_Kernel21_Valid_Out, channel58_Kernel21_Valid_Out, channel59_Kernel21_Valid_Out, channel60_Kernel21_Valid_Out, channel61_Kernel21_Valid_Out, channel62_Kernel21_Valid_Out, channel63_Kernel21_Valid_Out, channel64_Kernel21_Valid_Out;

	assign add_kernel21=channel1_Kernel21_Valid_Out & channel2_Kernel21_Valid_Out & channel3_Kernel21_Valid_Out & channel4_Kernel21_Valid_Out & channel5_Kernel21_Valid_Out & channel6_Kernel21_Valid_Out & channel7_Kernel21_Valid_Out & channel8_Kernel21_Valid_Out & channel9_Kernel21_Valid_Out & channel10_Kernel21_Valid_Out & channel11_Kernel21_Valid_Out & channel12_Kernel21_Valid_Out & channel13_Kernel21_Valid_Out & channel14_Kernel21_Valid_Out & channel15_Kernel21_Valid_Out & channel16_Kernel21_Valid_Out & channel17_Kernel21_Valid_Out & channel18_Kernel21_Valid_Out & channel19_Kernel21_Valid_Out & channel20_Kernel21_Valid_Out & channel21_Kernel21_Valid_Out & channel22_Kernel21_Valid_Out & channel23_Kernel21_Valid_Out & channel24_Kernel21_Valid_Out & channel25_Kernel21_Valid_Out & channel26_Kernel21_Valid_Out & channel27_Kernel21_Valid_Out & channel28_Kernel21_Valid_Out & channel29_Kernel21_Valid_Out & channel30_Kernel21_Valid_Out & channel31_Kernel21_Valid_Out & channel32_Kernel21_Valid_Out & channel33_Kernel21_Valid_Out & channel34_Kernel21_Valid_Out & channel35_Kernel21_Valid_Out & channel36_Kernel21_Valid_Out & channel37_Kernel21_Valid_Out & channel38_Kernel21_Valid_Out & channel39_Kernel21_Valid_Out & channel40_Kernel21_Valid_Out & channel41_Kernel21_Valid_Out & channel42_Kernel21_Valid_Out & channel43_Kernel21_Valid_Out & channel44_Kernel21_Valid_Out & channel45_Kernel21_Valid_Out & channel46_Kernel21_Valid_Out & channel47_Kernel21_Valid_Out & channel48_Kernel21_Valid_Out & channel49_Kernel21_Valid_Out & channel50_Kernel21_Valid_Out & channel51_Kernel21_Valid_Out & channel52_Kernel21_Valid_Out & channel53_Kernel21_Valid_Out & channel54_Kernel21_Valid_Out & channel55_Kernel21_Valid_Out & channel56_Kernel21_Valid_Out & channel57_Kernel21_Valid_Out & channel58_Kernel21_Valid_Out & channel59_Kernel21_Valid_Out & channel60_Kernel21_Valid_Out & channel61_Kernel21_Valid_Out & channel62_Kernel21_Valid_Out & channel63_Kernel21_Valid_Out & channel64_Kernel21_Valid_Out;

	wire channel1_Kernel22_Valid_Out, channel2_Kernel22_Valid_Out, channel3_Kernel22_Valid_Out, channel4_Kernel22_Valid_Out, channel5_Kernel22_Valid_Out, channel6_Kernel22_Valid_Out, channel7_Kernel22_Valid_Out, channel8_Kernel22_Valid_Out, channel9_Kernel22_Valid_Out, channel10_Kernel22_Valid_Out, channel11_Kernel22_Valid_Out, channel12_Kernel22_Valid_Out, channel13_Kernel22_Valid_Out, channel14_Kernel22_Valid_Out, channel15_Kernel22_Valid_Out, channel16_Kernel22_Valid_Out, channel17_Kernel22_Valid_Out, channel18_Kernel22_Valid_Out, channel19_Kernel22_Valid_Out, channel20_Kernel22_Valid_Out, channel21_Kernel22_Valid_Out, channel22_Kernel22_Valid_Out, channel23_Kernel22_Valid_Out, channel24_Kernel22_Valid_Out, channel25_Kernel22_Valid_Out, channel26_Kernel22_Valid_Out, channel27_Kernel22_Valid_Out, channel28_Kernel22_Valid_Out, channel29_Kernel22_Valid_Out, channel30_Kernel22_Valid_Out, channel31_Kernel22_Valid_Out, channel32_Kernel22_Valid_Out, channel33_Kernel22_Valid_Out, channel34_Kernel22_Valid_Out, channel35_Kernel22_Valid_Out, channel36_Kernel22_Valid_Out, channel37_Kernel22_Valid_Out, channel38_Kernel22_Valid_Out, channel39_Kernel22_Valid_Out, channel40_Kernel22_Valid_Out, channel41_Kernel22_Valid_Out, channel42_Kernel22_Valid_Out, channel43_Kernel22_Valid_Out, channel44_Kernel22_Valid_Out, channel45_Kernel22_Valid_Out, channel46_Kernel22_Valid_Out, channel47_Kernel22_Valid_Out, channel48_Kernel22_Valid_Out, channel49_Kernel22_Valid_Out, channel50_Kernel22_Valid_Out, channel51_Kernel22_Valid_Out, channel52_Kernel22_Valid_Out, channel53_Kernel22_Valid_Out, channel54_Kernel22_Valid_Out, channel55_Kernel22_Valid_Out, channel56_Kernel22_Valid_Out, channel57_Kernel22_Valid_Out, channel58_Kernel22_Valid_Out, channel59_Kernel22_Valid_Out, channel60_Kernel22_Valid_Out, channel61_Kernel22_Valid_Out, channel62_Kernel22_Valid_Out, channel63_Kernel22_Valid_Out, channel64_Kernel22_Valid_Out;

	assign add_kernel22=channel1_Kernel22_Valid_Out & channel2_Kernel22_Valid_Out & channel3_Kernel22_Valid_Out & channel4_Kernel22_Valid_Out & channel5_Kernel22_Valid_Out & channel6_Kernel22_Valid_Out & channel7_Kernel22_Valid_Out & channel8_Kernel22_Valid_Out & channel9_Kernel22_Valid_Out & channel10_Kernel22_Valid_Out & channel11_Kernel22_Valid_Out & channel12_Kernel22_Valid_Out & channel13_Kernel22_Valid_Out & channel14_Kernel22_Valid_Out & channel15_Kernel22_Valid_Out & channel16_Kernel22_Valid_Out & channel17_Kernel22_Valid_Out & channel18_Kernel22_Valid_Out & channel19_Kernel22_Valid_Out & channel20_Kernel22_Valid_Out & channel21_Kernel22_Valid_Out & channel22_Kernel22_Valid_Out & channel23_Kernel22_Valid_Out & channel24_Kernel22_Valid_Out & channel25_Kernel22_Valid_Out & channel26_Kernel22_Valid_Out & channel27_Kernel22_Valid_Out & channel28_Kernel22_Valid_Out & channel29_Kernel22_Valid_Out & channel30_Kernel22_Valid_Out & channel31_Kernel22_Valid_Out & channel32_Kernel22_Valid_Out & channel33_Kernel22_Valid_Out & channel34_Kernel22_Valid_Out & channel35_Kernel22_Valid_Out & channel36_Kernel22_Valid_Out & channel37_Kernel22_Valid_Out & channel38_Kernel22_Valid_Out & channel39_Kernel22_Valid_Out & channel40_Kernel22_Valid_Out & channel41_Kernel22_Valid_Out & channel42_Kernel22_Valid_Out & channel43_Kernel22_Valid_Out & channel44_Kernel22_Valid_Out & channel45_Kernel22_Valid_Out & channel46_Kernel22_Valid_Out & channel47_Kernel22_Valid_Out & channel48_Kernel22_Valid_Out & channel49_Kernel22_Valid_Out & channel50_Kernel22_Valid_Out & channel51_Kernel22_Valid_Out & channel52_Kernel22_Valid_Out & channel53_Kernel22_Valid_Out & channel54_Kernel22_Valid_Out & channel55_Kernel22_Valid_Out & channel56_Kernel22_Valid_Out & channel57_Kernel22_Valid_Out & channel58_Kernel22_Valid_Out & channel59_Kernel22_Valid_Out & channel60_Kernel22_Valid_Out & channel61_Kernel22_Valid_Out & channel62_Kernel22_Valid_Out & channel63_Kernel22_Valid_Out & channel64_Kernel22_Valid_Out;

	wire channel1_Kernel23_Valid_Out, channel2_Kernel23_Valid_Out, channel3_Kernel23_Valid_Out, channel4_Kernel23_Valid_Out, channel5_Kernel23_Valid_Out, channel6_Kernel23_Valid_Out, channel7_Kernel23_Valid_Out, channel8_Kernel23_Valid_Out, channel9_Kernel23_Valid_Out, channel10_Kernel23_Valid_Out, channel11_Kernel23_Valid_Out, channel12_Kernel23_Valid_Out, channel13_Kernel23_Valid_Out, channel14_Kernel23_Valid_Out, channel15_Kernel23_Valid_Out, channel16_Kernel23_Valid_Out, channel17_Kernel23_Valid_Out, channel18_Kernel23_Valid_Out, channel19_Kernel23_Valid_Out, channel20_Kernel23_Valid_Out, channel21_Kernel23_Valid_Out, channel22_Kernel23_Valid_Out, channel23_Kernel23_Valid_Out, channel24_Kernel23_Valid_Out, channel25_Kernel23_Valid_Out, channel26_Kernel23_Valid_Out, channel27_Kernel23_Valid_Out, channel28_Kernel23_Valid_Out, channel29_Kernel23_Valid_Out, channel30_Kernel23_Valid_Out, channel31_Kernel23_Valid_Out, channel32_Kernel23_Valid_Out, channel33_Kernel23_Valid_Out, channel34_Kernel23_Valid_Out, channel35_Kernel23_Valid_Out, channel36_Kernel23_Valid_Out, channel37_Kernel23_Valid_Out, channel38_Kernel23_Valid_Out, channel39_Kernel23_Valid_Out, channel40_Kernel23_Valid_Out, channel41_Kernel23_Valid_Out, channel42_Kernel23_Valid_Out, channel43_Kernel23_Valid_Out, channel44_Kernel23_Valid_Out, channel45_Kernel23_Valid_Out, channel46_Kernel23_Valid_Out, channel47_Kernel23_Valid_Out, channel48_Kernel23_Valid_Out, channel49_Kernel23_Valid_Out, channel50_Kernel23_Valid_Out, channel51_Kernel23_Valid_Out, channel52_Kernel23_Valid_Out, channel53_Kernel23_Valid_Out, channel54_Kernel23_Valid_Out, channel55_Kernel23_Valid_Out, channel56_Kernel23_Valid_Out, channel57_Kernel23_Valid_Out, channel58_Kernel23_Valid_Out, channel59_Kernel23_Valid_Out, channel60_Kernel23_Valid_Out, channel61_Kernel23_Valid_Out, channel62_Kernel23_Valid_Out, channel63_Kernel23_Valid_Out, channel64_Kernel23_Valid_Out;

	assign add_kernel23=channel1_Kernel23_Valid_Out & channel2_Kernel23_Valid_Out & channel3_Kernel23_Valid_Out & channel4_Kernel23_Valid_Out & channel5_Kernel23_Valid_Out & channel6_Kernel23_Valid_Out & channel7_Kernel23_Valid_Out & channel8_Kernel23_Valid_Out & channel9_Kernel23_Valid_Out & channel10_Kernel23_Valid_Out & channel11_Kernel23_Valid_Out & channel12_Kernel23_Valid_Out & channel13_Kernel23_Valid_Out & channel14_Kernel23_Valid_Out & channel15_Kernel23_Valid_Out & channel16_Kernel23_Valid_Out & channel17_Kernel23_Valid_Out & channel18_Kernel23_Valid_Out & channel19_Kernel23_Valid_Out & channel20_Kernel23_Valid_Out & channel21_Kernel23_Valid_Out & channel22_Kernel23_Valid_Out & channel23_Kernel23_Valid_Out & channel24_Kernel23_Valid_Out & channel25_Kernel23_Valid_Out & channel26_Kernel23_Valid_Out & channel27_Kernel23_Valid_Out & channel28_Kernel23_Valid_Out & channel29_Kernel23_Valid_Out & channel30_Kernel23_Valid_Out & channel31_Kernel23_Valid_Out & channel32_Kernel23_Valid_Out & channel33_Kernel23_Valid_Out & channel34_Kernel23_Valid_Out & channel35_Kernel23_Valid_Out & channel36_Kernel23_Valid_Out & channel37_Kernel23_Valid_Out & channel38_Kernel23_Valid_Out & channel39_Kernel23_Valid_Out & channel40_Kernel23_Valid_Out & channel41_Kernel23_Valid_Out & channel42_Kernel23_Valid_Out & channel43_Kernel23_Valid_Out & channel44_Kernel23_Valid_Out & channel45_Kernel23_Valid_Out & channel46_Kernel23_Valid_Out & channel47_Kernel23_Valid_Out & channel48_Kernel23_Valid_Out & channel49_Kernel23_Valid_Out & channel50_Kernel23_Valid_Out & channel51_Kernel23_Valid_Out & channel52_Kernel23_Valid_Out & channel53_Kernel23_Valid_Out & channel54_Kernel23_Valid_Out & channel55_Kernel23_Valid_Out & channel56_Kernel23_Valid_Out & channel57_Kernel23_Valid_Out & channel58_Kernel23_Valid_Out & channel59_Kernel23_Valid_Out & channel60_Kernel23_Valid_Out & channel61_Kernel23_Valid_Out & channel62_Kernel23_Valid_Out & channel63_Kernel23_Valid_Out & channel64_Kernel23_Valid_Out;

	wire channel1_Kernel24_Valid_Out, channel2_Kernel24_Valid_Out, channel3_Kernel24_Valid_Out, channel4_Kernel24_Valid_Out, channel5_Kernel24_Valid_Out, channel6_Kernel24_Valid_Out, channel7_Kernel24_Valid_Out, channel8_Kernel24_Valid_Out, channel9_Kernel24_Valid_Out, channel10_Kernel24_Valid_Out, channel11_Kernel24_Valid_Out, channel12_Kernel24_Valid_Out, channel13_Kernel24_Valid_Out, channel14_Kernel24_Valid_Out, channel15_Kernel24_Valid_Out, channel16_Kernel24_Valid_Out, channel17_Kernel24_Valid_Out, channel18_Kernel24_Valid_Out, channel19_Kernel24_Valid_Out, channel20_Kernel24_Valid_Out, channel21_Kernel24_Valid_Out, channel22_Kernel24_Valid_Out, channel23_Kernel24_Valid_Out, channel24_Kernel24_Valid_Out, channel25_Kernel24_Valid_Out, channel26_Kernel24_Valid_Out, channel27_Kernel24_Valid_Out, channel28_Kernel24_Valid_Out, channel29_Kernel24_Valid_Out, channel30_Kernel24_Valid_Out, channel31_Kernel24_Valid_Out, channel32_Kernel24_Valid_Out, channel33_Kernel24_Valid_Out, channel34_Kernel24_Valid_Out, channel35_Kernel24_Valid_Out, channel36_Kernel24_Valid_Out, channel37_Kernel24_Valid_Out, channel38_Kernel24_Valid_Out, channel39_Kernel24_Valid_Out, channel40_Kernel24_Valid_Out, channel41_Kernel24_Valid_Out, channel42_Kernel24_Valid_Out, channel43_Kernel24_Valid_Out, channel44_Kernel24_Valid_Out, channel45_Kernel24_Valid_Out, channel46_Kernel24_Valid_Out, channel47_Kernel24_Valid_Out, channel48_Kernel24_Valid_Out, channel49_Kernel24_Valid_Out, channel50_Kernel24_Valid_Out, channel51_Kernel24_Valid_Out, channel52_Kernel24_Valid_Out, channel53_Kernel24_Valid_Out, channel54_Kernel24_Valid_Out, channel55_Kernel24_Valid_Out, channel56_Kernel24_Valid_Out, channel57_Kernel24_Valid_Out, channel58_Kernel24_Valid_Out, channel59_Kernel24_Valid_Out, channel60_Kernel24_Valid_Out, channel61_Kernel24_Valid_Out, channel62_Kernel24_Valid_Out, channel63_Kernel24_Valid_Out, channel64_Kernel24_Valid_Out;

	assign add_kernel24=channel1_Kernel24_Valid_Out & channel2_Kernel24_Valid_Out & channel3_Kernel24_Valid_Out & channel4_Kernel24_Valid_Out & channel5_Kernel24_Valid_Out & channel6_Kernel24_Valid_Out & channel7_Kernel24_Valid_Out & channel8_Kernel24_Valid_Out & channel9_Kernel24_Valid_Out & channel10_Kernel24_Valid_Out & channel11_Kernel24_Valid_Out & channel12_Kernel24_Valid_Out & channel13_Kernel24_Valid_Out & channel14_Kernel24_Valid_Out & channel15_Kernel24_Valid_Out & channel16_Kernel24_Valid_Out & channel17_Kernel24_Valid_Out & channel18_Kernel24_Valid_Out & channel19_Kernel24_Valid_Out & channel20_Kernel24_Valid_Out & channel21_Kernel24_Valid_Out & channel22_Kernel24_Valid_Out & channel23_Kernel24_Valid_Out & channel24_Kernel24_Valid_Out & channel25_Kernel24_Valid_Out & channel26_Kernel24_Valid_Out & channel27_Kernel24_Valid_Out & channel28_Kernel24_Valid_Out & channel29_Kernel24_Valid_Out & channel30_Kernel24_Valid_Out & channel31_Kernel24_Valid_Out & channel32_Kernel24_Valid_Out & channel33_Kernel24_Valid_Out & channel34_Kernel24_Valid_Out & channel35_Kernel24_Valid_Out & channel36_Kernel24_Valid_Out & channel37_Kernel24_Valid_Out & channel38_Kernel24_Valid_Out & channel39_Kernel24_Valid_Out & channel40_Kernel24_Valid_Out & channel41_Kernel24_Valid_Out & channel42_Kernel24_Valid_Out & channel43_Kernel24_Valid_Out & channel44_Kernel24_Valid_Out & channel45_Kernel24_Valid_Out & channel46_Kernel24_Valid_Out & channel47_Kernel24_Valid_Out & channel48_Kernel24_Valid_Out & channel49_Kernel24_Valid_Out & channel50_Kernel24_Valid_Out & channel51_Kernel24_Valid_Out & channel52_Kernel24_Valid_Out & channel53_Kernel24_Valid_Out & channel54_Kernel24_Valid_Out & channel55_Kernel24_Valid_Out & channel56_Kernel24_Valid_Out & channel57_Kernel24_Valid_Out & channel58_Kernel24_Valid_Out & channel59_Kernel24_Valid_Out & channel60_Kernel24_Valid_Out & channel61_Kernel24_Valid_Out & channel62_Kernel24_Valid_Out & channel63_Kernel24_Valid_Out & channel64_Kernel24_Valid_Out;

	wire channel1_Kernel25_Valid_Out, channel2_Kernel25_Valid_Out, channel3_Kernel25_Valid_Out, channel4_Kernel25_Valid_Out, channel5_Kernel25_Valid_Out, channel6_Kernel25_Valid_Out, channel7_Kernel25_Valid_Out, channel8_Kernel25_Valid_Out, channel9_Kernel25_Valid_Out, channel10_Kernel25_Valid_Out, channel11_Kernel25_Valid_Out, channel12_Kernel25_Valid_Out, channel13_Kernel25_Valid_Out, channel14_Kernel25_Valid_Out, channel15_Kernel25_Valid_Out, channel16_Kernel25_Valid_Out, channel17_Kernel25_Valid_Out, channel18_Kernel25_Valid_Out, channel19_Kernel25_Valid_Out, channel20_Kernel25_Valid_Out, channel21_Kernel25_Valid_Out, channel22_Kernel25_Valid_Out, channel23_Kernel25_Valid_Out, channel24_Kernel25_Valid_Out, channel25_Kernel25_Valid_Out, channel26_Kernel25_Valid_Out, channel27_Kernel25_Valid_Out, channel28_Kernel25_Valid_Out, channel29_Kernel25_Valid_Out, channel30_Kernel25_Valid_Out, channel31_Kernel25_Valid_Out, channel32_Kernel25_Valid_Out, channel33_Kernel25_Valid_Out, channel34_Kernel25_Valid_Out, channel35_Kernel25_Valid_Out, channel36_Kernel25_Valid_Out, channel37_Kernel25_Valid_Out, channel38_Kernel25_Valid_Out, channel39_Kernel25_Valid_Out, channel40_Kernel25_Valid_Out, channel41_Kernel25_Valid_Out, channel42_Kernel25_Valid_Out, channel43_Kernel25_Valid_Out, channel44_Kernel25_Valid_Out, channel45_Kernel25_Valid_Out, channel46_Kernel25_Valid_Out, channel47_Kernel25_Valid_Out, channel48_Kernel25_Valid_Out, channel49_Kernel25_Valid_Out, channel50_Kernel25_Valid_Out, channel51_Kernel25_Valid_Out, channel52_Kernel25_Valid_Out, channel53_Kernel25_Valid_Out, channel54_Kernel25_Valid_Out, channel55_Kernel25_Valid_Out, channel56_Kernel25_Valid_Out, channel57_Kernel25_Valid_Out, channel58_Kernel25_Valid_Out, channel59_Kernel25_Valid_Out, channel60_Kernel25_Valid_Out, channel61_Kernel25_Valid_Out, channel62_Kernel25_Valid_Out, channel63_Kernel25_Valid_Out, channel64_Kernel25_Valid_Out;

	assign add_kernel25=channel1_Kernel25_Valid_Out & channel2_Kernel25_Valid_Out & channel3_Kernel25_Valid_Out & channel4_Kernel25_Valid_Out & channel5_Kernel25_Valid_Out & channel6_Kernel25_Valid_Out & channel7_Kernel25_Valid_Out & channel8_Kernel25_Valid_Out & channel9_Kernel25_Valid_Out & channel10_Kernel25_Valid_Out & channel11_Kernel25_Valid_Out & channel12_Kernel25_Valid_Out & channel13_Kernel25_Valid_Out & channel14_Kernel25_Valid_Out & channel15_Kernel25_Valid_Out & channel16_Kernel25_Valid_Out & channel17_Kernel25_Valid_Out & channel18_Kernel25_Valid_Out & channel19_Kernel25_Valid_Out & channel20_Kernel25_Valid_Out & channel21_Kernel25_Valid_Out & channel22_Kernel25_Valid_Out & channel23_Kernel25_Valid_Out & channel24_Kernel25_Valid_Out & channel25_Kernel25_Valid_Out & channel26_Kernel25_Valid_Out & channel27_Kernel25_Valid_Out & channel28_Kernel25_Valid_Out & channel29_Kernel25_Valid_Out & channel30_Kernel25_Valid_Out & channel31_Kernel25_Valid_Out & channel32_Kernel25_Valid_Out & channel33_Kernel25_Valid_Out & channel34_Kernel25_Valid_Out & channel35_Kernel25_Valid_Out & channel36_Kernel25_Valid_Out & channel37_Kernel25_Valid_Out & channel38_Kernel25_Valid_Out & channel39_Kernel25_Valid_Out & channel40_Kernel25_Valid_Out & channel41_Kernel25_Valid_Out & channel42_Kernel25_Valid_Out & channel43_Kernel25_Valid_Out & channel44_Kernel25_Valid_Out & channel45_Kernel25_Valid_Out & channel46_Kernel25_Valid_Out & channel47_Kernel25_Valid_Out & channel48_Kernel25_Valid_Out & channel49_Kernel25_Valid_Out & channel50_Kernel25_Valid_Out & channel51_Kernel25_Valid_Out & channel52_Kernel25_Valid_Out & channel53_Kernel25_Valid_Out & channel54_Kernel25_Valid_Out & channel55_Kernel25_Valid_Out & channel56_Kernel25_Valid_Out & channel57_Kernel25_Valid_Out & channel58_Kernel25_Valid_Out & channel59_Kernel25_Valid_Out & channel60_Kernel25_Valid_Out & channel61_Kernel25_Valid_Out & channel62_Kernel25_Valid_Out & channel63_Kernel25_Valid_Out & channel64_Kernel25_Valid_Out;

	wire channel1_Kernel26_Valid_Out, channel2_Kernel26_Valid_Out, channel3_Kernel26_Valid_Out, channel4_Kernel26_Valid_Out, channel5_Kernel26_Valid_Out, channel6_Kernel26_Valid_Out, channel7_Kernel26_Valid_Out, channel8_Kernel26_Valid_Out, channel9_Kernel26_Valid_Out, channel10_Kernel26_Valid_Out, channel11_Kernel26_Valid_Out, channel12_Kernel26_Valid_Out, channel13_Kernel26_Valid_Out, channel14_Kernel26_Valid_Out, channel15_Kernel26_Valid_Out, channel16_Kernel26_Valid_Out, channel17_Kernel26_Valid_Out, channel18_Kernel26_Valid_Out, channel19_Kernel26_Valid_Out, channel20_Kernel26_Valid_Out, channel21_Kernel26_Valid_Out, channel22_Kernel26_Valid_Out, channel23_Kernel26_Valid_Out, channel24_Kernel26_Valid_Out, channel25_Kernel26_Valid_Out, channel26_Kernel26_Valid_Out, channel27_Kernel26_Valid_Out, channel28_Kernel26_Valid_Out, channel29_Kernel26_Valid_Out, channel30_Kernel26_Valid_Out, channel31_Kernel26_Valid_Out, channel32_Kernel26_Valid_Out, channel33_Kernel26_Valid_Out, channel34_Kernel26_Valid_Out, channel35_Kernel26_Valid_Out, channel36_Kernel26_Valid_Out, channel37_Kernel26_Valid_Out, channel38_Kernel26_Valid_Out, channel39_Kernel26_Valid_Out, channel40_Kernel26_Valid_Out, channel41_Kernel26_Valid_Out, channel42_Kernel26_Valid_Out, channel43_Kernel26_Valid_Out, channel44_Kernel26_Valid_Out, channel45_Kernel26_Valid_Out, channel46_Kernel26_Valid_Out, channel47_Kernel26_Valid_Out, channel48_Kernel26_Valid_Out, channel49_Kernel26_Valid_Out, channel50_Kernel26_Valid_Out, channel51_Kernel26_Valid_Out, channel52_Kernel26_Valid_Out, channel53_Kernel26_Valid_Out, channel54_Kernel26_Valid_Out, channel55_Kernel26_Valid_Out, channel56_Kernel26_Valid_Out, channel57_Kernel26_Valid_Out, channel58_Kernel26_Valid_Out, channel59_Kernel26_Valid_Out, channel60_Kernel26_Valid_Out, channel61_Kernel26_Valid_Out, channel62_Kernel26_Valid_Out, channel63_Kernel26_Valid_Out, channel64_Kernel26_Valid_Out;

	assign add_kernel26=channel1_Kernel26_Valid_Out & channel2_Kernel26_Valid_Out & channel3_Kernel26_Valid_Out & channel4_Kernel26_Valid_Out & channel5_Kernel26_Valid_Out & channel6_Kernel26_Valid_Out & channel7_Kernel26_Valid_Out & channel8_Kernel26_Valid_Out & channel9_Kernel26_Valid_Out & channel10_Kernel26_Valid_Out & channel11_Kernel26_Valid_Out & channel12_Kernel26_Valid_Out & channel13_Kernel26_Valid_Out & channel14_Kernel26_Valid_Out & channel15_Kernel26_Valid_Out & channel16_Kernel26_Valid_Out & channel17_Kernel26_Valid_Out & channel18_Kernel26_Valid_Out & channel19_Kernel26_Valid_Out & channel20_Kernel26_Valid_Out & channel21_Kernel26_Valid_Out & channel22_Kernel26_Valid_Out & channel23_Kernel26_Valid_Out & channel24_Kernel26_Valid_Out & channel25_Kernel26_Valid_Out & channel26_Kernel26_Valid_Out & channel27_Kernel26_Valid_Out & channel28_Kernel26_Valid_Out & channel29_Kernel26_Valid_Out & channel30_Kernel26_Valid_Out & channel31_Kernel26_Valid_Out & channel32_Kernel26_Valid_Out & channel33_Kernel26_Valid_Out & channel34_Kernel26_Valid_Out & channel35_Kernel26_Valid_Out & channel36_Kernel26_Valid_Out & channel37_Kernel26_Valid_Out & channel38_Kernel26_Valid_Out & channel39_Kernel26_Valid_Out & channel40_Kernel26_Valid_Out & channel41_Kernel26_Valid_Out & channel42_Kernel26_Valid_Out & channel43_Kernel26_Valid_Out & channel44_Kernel26_Valid_Out & channel45_Kernel26_Valid_Out & channel46_Kernel26_Valid_Out & channel47_Kernel26_Valid_Out & channel48_Kernel26_Valid_Out & channel49_Kernel26_Valid_Out & channel50_Kernel26_Valid_Out & channel51_Kernel26_Valid_Out & channel52_Kernel26_Valid_Out & channel53_Kernel26_Valid_Out & channel54_Kernel26_Valid_Out & channel55_Kernel26_Valid_Out & channel56_Kernel26_Valid_Out & channel57_Kernel26_Valid_Out & channel58_Kernel26_Valid_Out & channel59_Kernel26_Valid_Out & channel60_Kernel26_Valid_Out & channel61_Kernel26_Valid_Out & channel62_Kernel26_Valid_Out & channel63_Kernel26_Valid_Out & channel64_Kernel26_Valid_Out;

	wire channel1_Kernel27_Valid_Out, channel2_Kernel27_Valid_Out, channel3_Kernel27_Valid_Out, channel4_Kernel27_Valid_Out, channel5_Kernel27_Valid_Out, channel6_Kernel27_Valid_Out, channel7_Kernel27_Valid_Out, channel8_Kernel27_Valid_Out, channel9_Kernel27_Valid_Out, channel10_Kernel27_Valid_Out, channel11_Kernel27_Valid_Out, channel12_Kernel27_Valid_Out, channel13_Kernel27_Valid_Out, channel14_Kernel27_Valid_Out, channel15_Kernel27_Valid_Out, channel16_Kernel27_Valid_Out, channel17_Kernel27_Valid_Out, channel18_Kernel27_Valid_Out, channel19_Kernel27_Valid_Out, channel20_Kernel27_Valid_Out, channel21_Kernel27_Valid_Out, channel22_Kernel27_Valid_Out, channel23_Kernel27_Valid_Out, channel24_Kernel27_Valid_Out, channel25_Kernel27_Valid_Out, channel26_Kernel27_Valid_Out, channel27_Kernel27_Valid_Out, channel28_Kernel27_Valid_Out, channel29_Kernel27_Valid_Out, channel30_Kernel27_Valid_Out, channel31_Kernel27_Valid_Out, channel32_Kernel27_Valid_Out, channel33_Kernel27_Valid_Out, channel34_Kernel27_Valid_Out, channel35_Kernel27_Valid_Out, channel36_Kernel27_Valid_Out, channel37_Kernel27_Valid_Out, channel38_Kernel27_Valid_Out, channel39_Kernel27_Valid_Out, channel40_Kernel27_Valid_Out, channel41_Kernel27_Valid_Out, channel42_Kernel27_Valid_Out, channel43_Kernel27_Valid_Out, channel44_Kernel27_Valid_Out, channel45_Kernel27_Valid_Out, channel46_Kernel27_Valid_Out, channel47_Kernel27_Valid_Out, channel48_Kernel27_Valid_Out, channel49_Kernel27_Valid_Out, channel50_Kernel27_Valid_Out, channel51_Kernel27_Valid_Out, channel52_Kernel27_Valid_Out, channel53_Kernel27_Valid_Out, channel54_Kernel27_Valid_Out, channel55_Kernel27_Valid_Out, channel56_Kernel27_Valid_Out, channel57_Kernel27_Valid_Out, channel58_Kernel27_Valid_Out, channel59_Kernel27_Valid_Out, channel60_Kernel27_Valid_Out, channel61_Kernel27_Valid_Out, channel62_Kernel27_Valid_Out, channel63_Kernel27_Valid_Out, channel64_Kernel27_Valid_Out;

	assign add_kernel27=channel1_Kernel27_Valid_Out & channel2_Kernel27_Valid_Out & channel3_Kernel27_Valid_Out & channel4_Kernel27_Valid_Out & channel5_Kernel27_Valid_Out & channel6_Kernel27_Valid_Out & channel7_Kernel27_Valid_Out & channel8_Kernel27_Valid_Out & channel9_Kernel27_Valid_Out & channel10_Kernel27_Valid_Out & channel11_Kernel27_Valid_Out & channel12_Kernel27_Valid_Out & channel13_Kernel27_Valid_Out & channel14_Kernel27_Valid_Out & channel15_Kernel27_Valid_Out & channel16_Kernel27_Valid_Out & channel17_Kernel27_Valid_Out & channel18_Kernel27_Valid_Out & channel19_Kernel27_Valid_Out & channel20_Kernel27_Valid_Out & channel21_Kernel27_Valid_Out & channel22_Kernel27_Valid_Out & channel23_Kernel27_Valid_Out & channel24_Kernel27_Valid_Out & channel25_Kernel27_Valid_Out & channel26_Kernel27_Valid_Out & channel27_Kernel27_Valid_Out & channel28_Kernel27_Valid_Out & channel29_Kernel27_Valid_Out & channel30_Kernel27_Valid_Out & channel31_Kernel27_Valid_Out & channel32_Kernel27_Valid_Out & channel33_Kernel27_Valid_Out & channel34_Kernel27_Valid_Out & channel35_Kernel27_Valid_Out & channel36_Kernel27_Valid_Out & channel37_Kernel27_Valid_Out & channel38_Kernel27_Valid_Out & channel39_Kernel27_Valid_Out & channel40_Kernel27_Valid_Out & channel41_Kernel27_Valid_Out & channel42_Kernel27_Valid_Out & channel43_Kernel27_Valid_Out & channel44_Kernel27_Valid_Out & channel45_Kernel27_Valid_Out & channel46_Kernel27_Valid_Out & channel47_Kernel27_Valid_Out & channel48_Kernel27_Valid_Out & channel49_Kernel27_Valid_Out & channel50_Kernel27_Valid_Out & channel51_Kernel27_Valid_Out & channel52_Kernel27_Valid_Out & channel53_Kernel27_Valid_Out & channel54_Kernel27_Valid_Out & channel55_Kernel27_Valid_Out & channel56_Kernel27_Valid_Out & channel57_Kernel27_Valid_Out & channel58_Kernel27_Valid_Out & channel59_Kernel27_Valid_Out & channel60_Kernel27_Valid_Out & channel61_Kernel27_Valid_Out & channel62_Kernel27_Valid_Out & channel63_Kernel27_Valid_Out & channel64_Kernel27_Valid_Out;

	wire channel1_Kernel28_Valid_Out, channel2_Kernel28_Valid_Out, channel3_Kernel28_Valid_Out, channel4_Kernel28_Valid_Out, channel5_Kernel28_Valid_Out, channel6_Kernel28_Valid_Out, channel7_Kernel28_Valid_Out, channel8_Kernel28_Valid_Out, channel9_Kernel28_Valid_Out, channel10_Kernel28_Valid_Out, channel11_Kernel28_Valid_Out, channel12_Kernel28_Valid_Out, channel13_Kernel28_Valid_Out, channel14_Kernel28_Valid_Out, channel15_Kernel28_Valid_Out, channel16_Kernel28_Valid_Out, channel17_Kernel28_Valid_Out, channel18_Kernel28_Valid_Out, channel19_Kernel28_Valid_Out, channel20_Kernel28_Valid_Out, channel21_Kernel28_Valid_Out, channel22_Kernel28_Valid_Out, channel23_Kernel28_Valid_Out, channel24_Kernel28_Valid_Out, channel25_Kernel28_Valid_Out, channel26_Kernel28_Valid_Out, channel27_Kernel28_Valid_Out, channel28_Kernel28_Valid_Out, channel29_Kernel28_Valid_Out, channel30_Kernel28_Valid_Out, channel31_Kernel28_Valid_Out, channel32_Kernel28_Valid_Out, channel33_Kernel28_Valid_Out, channel34_Kernel28_Valid_Out, channel35_Kernel28_Valid_Out, channel36_Kernel28_Valid_Out, channel37_Kernel28_Valid_Out, channel38_Kernel28_Valid_Out, channel39_Kernel28_Valid_Out, channel40_Kernel28_Valid_Out, channel41_Kernel28_Valid_Out, channel42_Kernel28_Valid_Out, channel43_Kernel28_Valid_Out, channel44_Kernel28_Valid_Out, channel45_Kernel28_Valid_Out, channel46_Kernel28_Valid_Out, channel47_Kernel28_Valid_Out, channel48_Kernel28_Valid_Out, channel49_Kernel28_Valid_Out, channel50_Kernel28_Valid_Out, channel51_Kernel28_Valid_Out, channel52_Kernel28_Valid_Out, channel53_Kernel28_Valid_Out, channel54_Kernel28_Valid_Out, channel55_Kernel28_Valid_Out, channel56_Kernel28_Valid_Out, channel57_Kernel28_Valid_Out, channel58_Kernel28_Valid_Out, channel59_Kernel28_Valid_Out, channel60_Kernel28_Valid_Out, channel61_Kernel28_Valid_Out, channel62_Kernel28_Valid_Out, channel63_Kernel28_Valid_Out, channel64_Kernel28_Valid_Out;

	assign add_kernel28=channel1_Kernel28_Valid_Out & channel2_Kernel28_Valid_Out & channel3_Kernel28_Valid_Out & channel4_Kernel28_Valid_Out & channel5_Kernel28_Valid_Out & channel6_Kernel28_Valid_Out & channel7_Kernel28_Valid_Out & channel8_Kernel28_Valid_Out & channel9_Kernel28_Valid_Out & channel10_Kernel28_Valid_Out & channel11_Kernel28_Valid_Out & channel12_Kernel28_Valid_Out & channel13_Kernel28_Valid_Out & channel14_Kernel28_Valid_Out & channel15_Kernel28_Valid_Out & channel16_Kernel28_Valid_Out & channel17_Kernel28_Valid_Out & channel18_Kernel28_Valid_Out & channel19_Kernel28_Valid_Out & channel20_Kernel28_Valid_Out & channel21_Kernel28_Valid_Out & channel22_Kernel28_Valid_Out & channel23_Kernel28_Valid_Out & channel24_Kernel28_Valid_Out & channel25_Kernel28_Valid_Out & channel26_Kernel28_Valid_Out & channel27_Kernel28_Valid_Out & channel28_Kernel28_Valid_Out & channel29_Kernel28_Valid_Out & channel30_Kernel28_Valid_Out & channel31_Kernel28_Valid_Out & channel32_Kernel28_Valid_Out & channel33_Kernel28_Valid_Out & channel34_Kernel28_Valid_Out & channel35_Kernel28_Valid_Out & channel36_Kernel28_Valid_Out & channel37_Kernel28_Valid_Out & channel38_Kernel28_Valid_Out & channel39_Kernel28_Valid_Out & channel40_Kernel28_Valid_Out & channel41_Kernel28_Valid_Out & channel42_Kernel28_Valid_Out & channel43_Kernel28_Valid_Out & channel44_Kernel28_Valid_Out & channel45_Kernel28_Valid_Out & channel46_Kernel28_Valid_Out & channel47_Kernel28_Valid_Out & channel48_Kernel28_Valid_Out & channel49_Kernel28_Valid_Out & channel50_Kernel28_Valid_Out & channel51_Kernel28_Valid_Out & channel52_Kernel28_Valid_Out & channel53_Kernel28_Valid_Out & channel54_Kernel28_Valid_Out & channel55_Kernel28_Valid_Out & channel56_Kernel28_Valid_Out & channel57_Kernel28_Valid_Out & channel58_Kernel28_Valid_Out & channel59_Kernel28_Valid_Out & channel60_Kernel28_Valid_Out & channel61_Kernel28_Valid_Out & channel62_Kernel28_Valid_Out & channel63_Kernel28_Valid_Out & channel64_Kernel28_Valid_Out;

	wire channel1_Kernel29_Valid_Out, channel2_Kernel29_Valid_Out, channel3_Kernel29_Valid_Out, channel4_Kernel29_Valid_Out, channel5_Kernel29_Valid_Out, channel6_Kernel29_Valid_Out, channel7_Kernel29_Valid_Out, channel8_Kernel29_Valid_Out, channel9_Kernel29_Valid_Out, channel10_Kernel29_Valid_Out, channel11_Kernel29_Valid_Out, channel12_Kernel29_Valid_Out, channel13_Kernel29_Valid_Out, channel14_Kernel29_Valid_Out, channel15_Kernel29_Valid_Out, channel16_Kernel29_Valid_Out, channel17_Kernel29_Valid_Out, channel18_Kernel29_Valid_Out, channel19_Kernel29_Valid_Out, channel20_Kernel29_Valid_Out, channel21_Kernel29_Valid_Out, channel22_Kernel29_Valid_Out, channel23_Kernel29_Valid_Out, channel24_Kernel29_Valid_Out, channel25_Kernel29_Valid_Out, channel26_Kernel29_Valid_Out, channel27_Kernel29_Valid_Out, channel28_Kernel29_Valid_Out, channel29_Kernel29_Valid_Out, channel30_Kernel29_Valid_Out, channel31_Kernel29_Valid_Out, channel32_Kernel29_Valid_Out, channel33_Kernel29_Valid_Out, channel34_Kernel29_Valid_Out, channel35_Kernel29_Valid_Out, channel36_Kernel29_Valid_Out, channel37_Kernel29_Valid_Out, channel38_Kernel29_Valid_Out, channel39_Kernel29_Valid_Out, channel40_Kernel29_Valid_Out, channel41_Kernel29_Valid_Out, channel42_Kernel29_Valid_Out, channel43_Kernel29_Valid_Out, channel44_Kernel29_Valid_Out, channel45_Kernel29_Valid_Out, channel46_Kernel29_Valid_Out, channel47_Kernel29_Valid_Out, channel48_Kernel29_Valid_Out, channel49_Kernel29_Valid_Out, channel50_Kernel29_Valid_Out, channel51_Kernel29_Valid_Out, channel52_Kernel29_Valid_Out, channel53_Kernel29_Valid_Out, channel54_Kernel29_Valid_Out, channel55_Kernel29_Valid_Out, channel56_Kernel29_Valid_Out, channel57_Kernel29_Valid_Out, channel58_Kernel29_Valid_Out, channel59_Kernel29_Valid_Out, channel60_Kernel29_Valid_Out, channel61_Kernel29_Valid_Out, channel62_Kernel29_Valid_Out, channel63_Kernel29_Valid_Out, channel64_Kernel29_Valid_Out;

	assign add_kernel29=channel1_Kernel29_Valid_Out & channel2_Kernel29_Valid_Out & channel3_Kernel29_Valid_Out & channel4_Kernel29_Valid_Out & channel5_Kernel29_Valid_Out & channel6_Kernel29_Valid_Out & channel7_Kernel29_Valid_Out & channel8_Kernel29_Valid_Out & channel9_Kernel29_Valid_Out & channel10_Kernel29_Valid_Out & channel11_Kernel29_Valid_Out & channel12_Kernel29_Valid_Out & channel13_Kernel29_Valid_Out & channel14_Kernel29_Valid_Out & channel15_Kernel29_Valid_Out & channel16_Kernel29_Valid_Out & channel17_Kernel29_Valid_Out & channel18_Kernel29_Valid_Out & channel19_Kernel29_Valid_Out & channel20_Kernel29_Valid_Out & channel21_Kernel29_Valid_Out & channel22_Kernel29_Valid_Out & channel23_Kernel29_Valid_Out & channel24_Kernel29_Valid_Out & channel25_Kernel29_Valid_Out & channel26_Kernel29_Valid_Out & channel27_Kernel29_Valid_Out & channel28_Kernel29_Valid_Out & channel29_Kernel29_Valid_Out & channel30_Kernel29_Valid_Out & channel31_Kernel29_Valid_Out & channel32_Kernel29_Valid_Out & channel33_Kernel29_Valid_Out & channel34_Kernel29_Valid_Out & channel35_Kernel29_Valid_Out & channel36_Kernel29_Valid_Out & channel37_Kernel29_Valid_Out & channel38_Kernel29_Valid_Out & channel39_Kernel29_Valid_Out & channel40_Kernel29_Valid_Out & channel41_Kernel29_Valid_Out & channel42_Kernel29_Valid_Out & channel43_Kernel29_Valid_Out & channel44_Kernel29_Valid_Out & channel45_Kernel29_Valid_Out & channel46_Kernel29_Valid_Out & channel47_Kernel29_Valid_Out & channel48_Kernel29_Valid_Out & channel49_Kernel29_Valid_Out & channel50_Kernel29_Valid_Out & channel51_Kernel29_Valid_Out & channel52_Kernel29_Valid_Out & channel53_Kernel29_Valid_Out & channel54_Kernel29_Valid_Out & channel55_Kernel29_Valid_Out & channel56_Kernel29_Valid_Out & channel57_Kernel29_Valid_Out & channel58_Kernel29_Valid_Out & channel59_Kernel29_Valid_Out & channel60_Kernel29_Valid_Out & channel61_Kernel29_Valid_Out & channel62_Kernel29_Valid_Out & channel63_Kernel29_Valid_Out & channel64_Kernel29_Valid_Out;

	wire channel1_Kernel30_Valid_Out, channel2_Kernel30_Valid_Out, channel3_Kernel30_Valid_Out, channel4_Kernel30_Valid_Out, channel5_Kernel30_Valid_Out, channel6_Kernel30_Valid_Out, channel7_Kernel30_Valid_Out, channel8_Kernel30_Valid_Out, channel9_Kernel30_Valid_Out, channel10_Kernel30_Valid_Out, channel11_Kernel30_Valid_Out, channel12_Kernel30_Valid_Out, channel13_Kernel30_Valid_Out, channel14_Kernel30_Valid_Out, channel15_Kernel30_Valid_Out, channel16_Kernel30_Valid_Out, channel17_Kernel30_Valid_Out, channel18_Kernel30_Valid_Out, channel19_Kernel30_Valid_Out, channel20_Kernel30_Valid_Out, channel21_Kernel30_Valid_Out, channel22_Kernel30_Valid_Out, channel23_Kernel30_Valid_Out, channel24_Kernel30_Valid_Out, channel25_Kernel30_Valid_Out, channel26_Kernel30_Valid_Out, channel27_Kernel30_Valid_Out, channel28_Kernel30_Valid_Out, channel29_Kernel30_Valid_Out, channel30_Kernel30_Valid_Out, channel31_Kernel30_Valid_Out, channel32_Kernel30_Valid_Out, channel33_Kernel30_Valid_Out, channel34_Kernel30_Valid_Out, channel35_Kernel30_Valid_Out, channel36_Kernel30_Valid_Out, channel37_Kernel30_Valid_Out, channel38_Kernel30_Valid_Out, channel39_Kernel30_Valid_Out, channel40_Kernel30_Valid_Out, channel41_Kernel30_Valid_Out, channel42_Kernel30_Valid_Out, channel43_Kernel30_Valid_Out, channel44_Kernel30_Valid_Out, channel45_Kernel30_Valid_Out, channel46_Kernel30_Valid_Out, channel47_Kernel30_Valid_Out, channel48_Kernel30_Valid_Out, channel49_Kernel30_Valid_Out, channel50_Kernel30_Valid_Out, channel51_Kernel30_Valid_Out, channel52_Kernel30_Valid_Out, channel53_Kernel30_Valid_Out, channel54_Kernel30_Valid_Out, channel55_Kernel30_Valid_Out, channel56_Kernel30_Valid_Out, channel57_Kernel30_Valid_Out, channel58_Kernel30_Valid_Out, channel59_Kernel30_Valid_Out, channel60_Kernel30_Valid_Out, channel61_Kernel30_Valid_Out, channel62_Kernel30_Valid_Out, channel63_Kernel30_Valid_Out, channel64_Kernel30_Valid_Out;

	assign add_kernel30=channel1_Kernel30_Valid_Out & channel2_Kernel30_Valid_Out & channel3_Kernel30_Valid_Out & channel4_Kernel30_Valid_Out & channel5_Kernel30_Valid_Out & channel6_Kernel30_Valid_Out & channel7_Kernel30_Valid_Out & channel8_Kernel30_Valid_Out & channel9_Kernel30_Valid_Out & channel10_Kernel30_Valid_Out & channel11_Kernel30_Valid_Out & channel12_Kernel30_Valid_Out & channel13_Kernel30_Valid_Out & channel14_Kernel30_Valid_Out & channel15_Kernel30_Valid_Out & channel16_Kernel30_Valid_Out & channel17_Kernel30_Valid_Out & channel18_Kernel30_Valid_Out & channel19_Kernel30_Valid_Out & channel20_Kernel30_Valid_Out & channel21_Kernel30_Valid_Out & channel22_Kernel30_Valid_Out & channel23_Kernel30_Valid_Out & channel24_Kernel30_Valid_Out & channel25_Kernel30_Valid_Out & channel26_Kernel30_Valid_Out & channel27_Kernel30_Valid_Out & channel28_Kernel30_Valid_Out & channel29_Kernel30_Valid_Out & channel30_Kernel30_Valid_Out & channel31_Kernel30_Valid_Out & channel32_Kernel30_Valid_Out & channel33_Kernel30_Valid_Out & channel34_Kernel30_Valid_Out & channel35_Kernel30_Valid_Out & channel36_Kernel30_Valid_Out & channel37_Kernel30_Valid_Out & channel38_Kernel30_Valid_Out & channel39_Kernel30_Valid_Out & channel40_Kernel30_Valid_Out & channel41_Kernel30_Valid_Out & channel42_Kernel30_Valid_Out & channel43_Kernel30_Valid_Out & channel44_Kernel30_Valid_Out & channel45_Kernel30_Valid_Out & channel46_Kernel30_Valid_Out & channel47_Kernel30_Valid_Out & channel48_Kernel30_Valid_Out & channel49_Kernel30_Valid_Out & channel50_Kernel30_Valid_Out & channel51_Kernel30_Valid_Out & channel52_Kernel30_Valid_Out & channel53_Kernel30_Valid_Out & channel54_Kernel30_Valid_Out & channel55_Kernel30_Valid_Out & channel56_Kernel30_Valid_Out & channel57_Kernel30_Valid_Out & channel58_Kernel30_Valid_Out & channel59_Kernel30_Valid_Out & channel60_Kernel30_Valid_Out & channel61_Kernel30_Valid_Out & channel62_Kernel30_Valid_Out & channel63_Kernel30_Valid_Out & channel64_Kernel30_Valid_Out;

	wire channel1_Kernel31_Valid_Out, channel2_Kernel31_Valid_Out, channel3_Kernel31_Valid_Out, channel4_Kernel31_Valid_Out, channel5_Kernel31_Valid_Out, channel6_Kernel31_Valid_Out, channel7_Kernel31_Valid_Out, channel8_Kernel31_Valid_Out, channel9_Kernel31_Valid_Out, channel10_Kernel31_Valid_Out, channel11_Kernel31_Valid_Out, channel12_Kernel31_Valid_Out, channel13_Kernel31_Valid_Out, channel14_Kernel31_Valid_Out, channel15_Kernel31_Valid_Out, channel16_Kernel31_Valid_Out, channel17_Kernel31_Valid_Out, channel18_Kernel31_Valid_Out, channel19_Kernel31_Valid_Out, channel20_Kernel31_Valid_Out, channel21_Kernel31_Valid_Out, channel22_Kernel31_Valid_Out, channel23_Kernel31_Valid_Out, channel24_Kernel31_Valid_Out, channel25_Kernel31_Valid_Out, channel26_Kernel31_Valid_Out, channel27_Kernel31_Valid_Out, channel28_Kernel31_Valid_Out, channel29_Kernel31_Valid_Out, channel30_Kernel31_Valid_Out, channel31_Kernel31_Valid_Out, channel32_Kernel31_Valid_Out, channel33_Kernel31_Valid_Out, channel34_Kernel31_Valid_Out, channel35_Kernel31_Valid_Out, channel36_Kernel31_Valid_Out, channel37_Kernel31_Valid_Out, channel38_Kernel31_Valid_Out, channel39_Kernel31_Valid_Out, channel40_Kernel31_Valid_Out, channel41_Kernel31_Valid_Out, channel42_Kernel31_Valid_Out, channel43_Kernel31_Valid_Out, channel44_Kernel31_Valid_Out, channel45_Kernel31_Valid_Out, channel46_Kernel31_Valid_Out, channel47_Kernel31_Valid_Out, channel48_Kernel31_Valid_Out, channel49_Kernel31_Valid_Out, channel50_Kernel31_Valid_Out, channel51_Kernel31_Valid_Out, channel52_Kernel31_Valid_Out, channel53_Kernel31_Valid_Out, channel54_Kernel31_Valid_Out, channel55_Kernel31_Valid_Out, channel56_Kernel31_Valid_Out, channel57_Kernel31_Valid_Out, channel58_Kernel31_Valid_Out, channel59_Kernel31_Valid_Out, channel60_Kernel31_Valid_Out, channel61_Kernel31_Valid_Out, channel62_Kernel31_Valid_Out, channel63_Kernel31_Valid_Out, channel64_Kernel31_Valid_Out;

	assign add_kernel31=channel1_Kernel31_Valid_Out & channel2_Kernel31_Valid_Out & channel3_Kernel31_Valid_Out & channel4_Kernel31_Valid_Out & channel5_Kernel31_Valid_Out & channel6_Kernel31_Valid_Out & channel7_Kernel31_Valid_Out & channel8_Kernel31_Valid_Out & channel9_Kernel31_Valid_Out & channel10_Kernel31_Valid_Out & channel11_Kernel31_Valid_Out & channel12_Kernel31_Valid_Out & channel13_Kernel31_Valid_Out & channel14_Kernel31_Valid_Out & channel15_Kernel31_Valid_Out & channel16_Kernel31_Valid_Out & channel17_Kernel31_Valid_Out & channel18_Kernel31_Valid_Out & channel19_Kernel31_Valid_Out & channel20_Kernel31_Valid_Out & channel21_Kernel31_Valid_Out & channel22_Kernel31_Valid_Out & channel23_Kernel31_Valid_Out & channel24_Kernel31_Valid_Out & channel25_Kernel31_Valid_Out & channel26_Kernel31_Valid_Out & channel27_Kernel31_Valid_Out & channel28_Kernel31_Valid_Out & channel29_Kernel31_Valid_Out & channel30_Kernel31_Valid_Out & channel31_Kernel31_Valid_Out & channel32_Kernel31_Valid_Out & channel33_Kernel31_Valid_Out & channel34_Kernel31_Valid_Out & channel35_Kernel31_Valid_Out & channel36_Kernel31_Valid_Out & channel37_Kernel31_Valid_Out & channel38_Kernel31_Valid_Out & channel39_Kernel31_Valid_Out & channel40_Kernel31_Valid_Out & channel41_Kernel31_Valid_Out & channel42_Kernel31_Valid_Out & channel43_Kernel31_Valid_Out & channel44_Kernel31_Valid_Out & channel45_Kernel31_Valid_Out & channel46_Kernel31_Valid_Out & channel47_Kernel31_Valid_Out & channel48_Kernel31_Valid_Out & channel49_Kernel31_Valid_Out & channel50_Kernel31_Valid_Out & channel51_Kernel31_Valid_Out & channel52_Kernel31_Valid_Out & channel53_Kernel31_Valid_Out & channel54_Kernel31_Valid_Out & channel55_Kernel31_Valid_Out & channel56_Kernel31_Valid_Out & channel57_Kernel31_Valid_Out & channel58_Kernel31_Valid_Out & channel59_Kernel31_Valid_Out & channel60_Kernel31_Valid_Out & channel61_Kernel31_Valid_Out & channel62_Kernel31_Valid_Out & channel63_Kernel31_Valid_Out & channel64_Kernel31_Valid_Out;

	wire channel1_Kernel32_Valid_Out, channel2_Kernel32_Valid_Out, channel3_Kernel32_Valid_Out, channel4_Kernel32_Valid_Out, channel5_Kernel32_Valid_Out, channel6_Kernel32_Valid_Out, channel7_Kernel32_Valid_Out, channel8_Kernel32_Valid_Out, channel9_Kernel32_Valid_Out, channel10_Kernel32_Valid_Out, channel11_Kernel32_Valid_Out, channel12_Kernel32_Valid_Out, channel13_Kernel32_Valid_Out, channel14_Kernel32_Valid_Out, channel15_Kernel32_Valid_Out, channel16_Kernel32_Valid_Out, channel17_Kernel32_Valid_Out, channel18_Kernel32_Valid_Out, channel19_Kernel32_Valid_Out, channel20_Kernel32_Valid_Out, channel21_Kernel32_Valid_Out, channel22_Kernel32_Valid_Out, channel23_Kernel32_Valid_Out, channel24_Kernel32_Valid_Out, channel25_Kernel32_Valid_Out, channel26_Kernel32_Valid_Out, channel27_Kernel32_Valid_Out, channel28_Kernel32_Valid_Out, channel29_Kernel32_Valid_Out, channel30_Kernel32_Valid_Out, channel31_Kernel32_Valid_Out, channel32_Kernel32_Valid_Out, channel33_Kernel32_Valid_Out, channel34_Kernel32_Valid_Out, channel35_Kernel32_Valid_Out, channel36_Kernel32_Valid_Out, channel37_Kernel32_Valid_Out, channel38_Kernel32_Valid_Out, channel39_Kernel32_Valid_Out, channel40_Kernel32_Valid_Out, channel41_Kernel32_Valid_Out, channel42_Kernel32_Valid_Out, channel43_Kernel32_Valid_Out, channel44_Kernel32_Valid_Out, channel45_Kernel32_Valid_Out, channel46_Kernel32_Valid_Out, channel47_Kernel32_Valid_Out, channel48_Kernel32_Valid_Out, channel49_Kernel32_Valid_Out, channel50_Kernel32_Valid_Out, channel51_Kernel32_Valid_Out, channel52_Kernel32_Valid_Out, channel53_Kernel32_Valid_Out, channel54_Kernel32_Valid_Out, channel55_Kernel32_Valid_Out, channel56_Kernel32_Valid_Out, channel57_Kernel32_Valid_Out, channel58_Kernel32_Valid_Out, channel59_Kernel32_Valid_Out, channel60_Kernel32_Valid_Out, channel61_Kernel32_Valid_Out, channel62_Kernel32_Valid_Out, channel63_Kernel32_Valid_Out, channel64_Kernel32_Valid_Out;

	assign add_kernel32=channel1_Kernel32_Valid_Out & channel2_Kernel32_Valid_Out & channel3_Kernel32_Valid_Out & channel4_Kernel32_Valid_Out & channel5_Kernel32_Valid_Out & channel6_Kernel32_Valid_Out & channel7_Kernel32_Valid_Out & channel8_Kernel32_Valid_Out & channel9_Kernel32_Valid_Out & channel10_Kernel32_Valid_Out & channel11_Kernel32_Valid_Out & channel12_Kernel32_Valid_Out & channel13_Kernel32_Valid_Out & channel14_Kernel32_Valid_Out & channel15_Kernel32_Valid_Out & channel16_Kernel32_Valid_Out & channel17_Kernel32_Valid_Out & channel18_Kernel32_Valid_Out & channel19_Kernel32_Valid_Out & channel20_Kernel32_Valid_Out & channel21_Kernel32_Valid_Out & channel22_Kernel32_Valid_Out & channel23_Kernel32_Valid_Out & channel24_Kernel32_Valid_Out & channel25_Kernel32_Valid_Out & channel26_Kernel32_Valid_Out & channel27_Kernel32_Valid_Out & channel28_Kernel32_Valid_Out & channel29_Kernel32_Valid_Out & channel30_Kernel32_Valid_Out & channel31_Kernel32_Valid_Out & channel32_Kernel32_Valid_Out & channel33_Kernel32_Valid_Out & channel34_Kernel32_Valid_Out & channel35_Kernel32_Valid_Out & channel36_Kernel32_Valid_Out & channel37_Kernel32_Valid_Out & channel38_Kernel32_Valid_Out & channel39_Kernel32_Valid_Out & channel40_Kernel32_Valid_Out & channel41_Kernel32_Valid_Out & channel42_Kernel32_Valid_Out & channel43_Kernel32_Valid_Out & channel44_Kernel32_Valid_Out & channel45_Kernel32_Valid_Out & channel46_Kernel32_Valid_Out & channel47_Kernel32_Valid_Out & channel48_Kernel32_Valid_Out & channel49_Kernel32_Valid_Out & channel50_Kernel32_Valid_Out & channel51_Kernel32_Valid_Out & channel52_Kernel32_Valid_Out & channel53_Kernel32_Valid_Out & channel54_Kernel32_Valid_Out & channel55_Kernel32_Valid_Out & channel56_Kernel32_Valid_Out & channel57_Kernel32_Valid_Out & channel58_Kernel32_Valid_Out & channel59_Kernel32_Valid_Out & channel60_Kernel32_Valid_Out & channel61_Kernel32_Valid_Out & channel62_Kernel32_Valid_Out & channel63_Kernel32_Valid_Out & channel64_Kernel32_Valid_Out;

	wire channel1_Kernel33_Valid_Out, channel2_Kernel33_Valid_Out, channel3_Kernel33_Valid_Out, channel4_Kernel33_Valid_Out, channel5_Kernel33_Valid_Out, channel6_Kernel33_Valid_Out, channel7_Kernel33_Valid_Out, channel8_Kernel33_Valid_Out, channel9_Kernel33_Valid_Out, channel10_Kernel33_Valid_Out, channel11_Kernel33_Valid_Out, channel12_Kernel33_Valid_Out, channel13_Kernel33_Valid_Out, channel14_Kernel33_Valid_Out, channel15_Kernel33_Valid_Out, channel16_Kernel33_Valid_Out, channel17_Kernel33_Valid_Out, channel18_Kernel33_Valid_Out, channel19_Kernel33_Valid_Out, channel20_Kernel33_Valid_Out, channel21_Kernel33_Valid_Out, channel22_Kernel33_Valid_Out, channel23_Kernel33_Valid_Out, channel24_Kernel33_Valid_Out, channel25_Kernel33_Valid_Out, channel26_Kernel33_Valid_Out, channel27_Kernel33_Valid_Out, channel28_Kernel33_Valid_Out, channel29_Kernel33_Valid_Out, channel30_Kernel33_Valid_Out, channel31_Kernel33_Valid_Out, channel32_Kernel33_Valid_Out, channel33_Kernel33_Valid_Out, channel34_Kernel33_Valid_Out, channel35_Kernel33_Valid_Out, channel36_Kernel33_Valid_Out, channel37_Kernel33_Valid_Out, channel38_Kernel33_Valid_Out, channel39_Kernel33_Valid_Out, channel40_Kernel33_Valid_Out, channel41_Kernel33_Valid_Out, channel42_Kernel33_Valid_Out, channel43_Kernel33_Valid_Out, channel44_Kernel33_Valid_Out, channel45_Kernel33_Valid_Out, channel46_Kernel33_Valid_Out, channel47_Kernel33_Valid_Out, channel48_Kernel33_Valid_Out, channel49_Kernel33_Valid_Out, channel50_Kernel33_Valid_Out, channel51_Kernel33_Valid_Out, channel52_Kernel33_Valid_Out, channel53_Kernel33_Valid_Out, channel54_Kernel33_Valid_Out, channel55_Kernel33_Valid_Out, channel56_Kernel33_Valid_Out, channel57_Kernel33_Valid_Out, channel58_Kernel33_Valid_Out, channel59_Kernel33_Valid_Out, channel60_Kernel33_Valid_Out, channel61_Kernel33_Valid_Out, channel62_Kernel33_Valid_Out, channel63_Kernel33_Valid_Out, channel64_Kernel33_Valid_Out;

	assign add_kernel33=channel1_Kernel33_Valid_Out & channel2_Kernel33_Valid_Out & channel3_Kernel33_Valid_Out & channel4_Kernel33_Valid_Out & channel5_Kernel33_Valid_Out & channel6_Kernel33_Valid_Out & channel7_Kernel33_Valid_Out & channel8_Kernel33_Valid_Out & channel9_Kernel33_Valid_Out & channel10_Kernel33_Valid_Out & channel11_Kernel33_Valid_Out & channel12_Kernel33_Valid_Out & channel13_Kernel33_Valid_Out & channel14_Kernel33_Valid_Out & channel15_Kernel33_Valid_Out & channel16_Kernel33_Valid_Out & channel17_Kernel33_Valid_Out & channel18_Kernel33_Valid_Out & channel19_Kernel33_Valid_Out & channel20_Kernel33_Valid_Out & channel21_Kernel33_Valid_Out & channel22_Kernel33_Valid_Out & channel23_Kernel33_Valid_Out & channel24_Kernel33_Valid_Out & channel25_Kernel33_Valid_Out & channel26_Kernel33_Valid_Out & channel27_Kernel33_Valid_Out & channel28_Kernel33_Valid_Out & channel29_Kernel33_Valid_Out & channel30_Kernel33_Valid_Out & channel31_Kernel33_Valid_Out & channel32_Kernel33_Valid_Out & channel33_Kernel33_Valid_Out & channel34_Kernel33_Valid_Out & channel35_Kernel33_Valid_Out & channel36_Kernel33_Valid_Out & channel37_Kernel33_Valid_Out & channel38_Kernel33_Valid_Out & channel39_Kernel33_Valid_Out & channel40_Kernel33_Valid_Out & channel41_Kernel33_Valid_Out & channel42_Kernel33_Valid_Out & channel43_Kernel33_Valid_Out & channel44_Kernel33_Valid_Out & channel45_Kernel33_Valid_Out & channel46_Kernel33_Valid_Out & channel47_Kernel33_Valid_Out & channel48_Kernel33_Valid_Out & channel49_Kernel33_Valid_Out & channel50_Kernel33_Valid_Out & channel51_Kernel33_Valid_Out & channel52_Kernel33_Valid_Out & channel53_Kernel33_Valid_Out & channel54_Kernel33_Valid_Out & channel55_Kernel33_Valid_Out & channel56_Kernel33_Valid_Out & channel57_Kernel33_Valid_Out & channel58_Kernel33_Valid_Out & channel59_Kernel33_Valid_Out & channel60_Kernel33_Valid_Out & channel61_Kernel33_Valid_Out & channel62_Kernel33_Valid_Out & channel63_Kernel33_Valid_Out & channel64_Kernel33_Valid_Out;

	wire channel1_Kernel34_Valid_Out, channel2_Kernel34_Valid_Out, channel3_Kernel34_Valid_Out, channel4_Kernel34_Valid_Out, channel5_Kernel34_Valid_Out, channel6_Kernel34_Valid_Out, channel7_Kernel34_Valid_Out, channel8_Kernel34_Valid_Out, channel9_Kernel34_Valid_Out, channel10_Kernel34_Valid_Out, channel11_Kernel34_Valid_Out, channel12_Kernel34_Valid_Out, channel13_Kernel34_Valid_Out, channel14_Kernel34_Valid_Out, channel15_Kernel34_Valid_Out, channel16_Kernel34_Valid_Out, channel17_Kernel34_Valid_Out, channel18_Kernel34_Valid_Out, channel19_Kernel34_Valid_Out, channel20_Kernel34_Valid_Out, channel21_Kernel34_Valid_Out, channel22_Kernel34_Valid_Out, channel23_Kernel34_Valid_Out, channel24_Kernel34_Valid_Out, channel25_Kernel34_Valid_Out, channel26_Kernel34_Valid_Out, channel27_Kernel34_Valid_Out, channel28_Kernel34_Valid_Out, channel29_Kernel34_Valid_Out, channel30_Kernel34_Valid_Out, channel31_Kernel34_Valid_Out, channel32_Kernel34_Valid_Out, channel33_Kernel34_Valid_Out, channel34_Kernel34_Valid_Out, channel35_Kernel34_Valid_Out, channel36_Kernel34_Valid_Out, channel37_Kernel34_Valid_Out, channel38_Kernel34_Valid_Out, channel39_Kernel34_Valid_Out, channel40_Kernel34_Valid_Out, channel41_Kernel34_Valid_Out, channel42_Kernel34_Valid_Out, channel43_Kernel34_Valid_Out, channel44_Kernel34_Valid_Out, channel45_Kernel34_Valid_Out, channel46_Kernel34_Valid_Out, channel47_Kernel34_Valid_Out, channel48_Kernel34_Valid_Out, channel49_Kernel34_Valid_Out, channel50_Kernel34_Valid_Out, channel51_Kernel34_Valid_Out, channel52_Kernel34_Valid_Out, channel53_Kernel34_Valid_Out, channel54_Kernel34_Valid_Out, channel55_Kernel34_Valid_Out, channel56_Kernel34_Valid_Out, channel57_Kernel34_Valid_Out, channel58_Kernel34_Valid_Out, channel59_Kernel34_Valid_Out, channel60_Kernel34_Valid_Out, channel61_Kernel34_Valid_Out, channel62_Kernel34_Valid_Out, channel63_Kernel34_Valid_Out, channel64_Kernel34_Valid_Out;

	assign add_kernel34=channel1_Kernel34_Valid_Out & channel2_Kernel34_Valid_Out & channel3_Kernel34_Valid_Out & channel4_Kernel34_Valid_Out & channel5_Kernel34_Valid_Out & channel6_Kernel34_Valid_Out & channel7_Kernel34_Valid_Out & channel8_Kernel34_Valid_Out & channel9_Kernel34_Valid_Out & channel10_Kernel34_Valid_Out & channel11_Kernel34_Valid_Out & channel12_Kernel34_Valid_Out & channel13_Kernel34_Valid_Out & channel14_Kernel34_Valid_Out & channel15_Kernel34_Valid_Out & channel16_Kernel34_Valid_Out & channel17_Kernel34_Valid_Out & channel18_Kernel34_Valid_Out & channel19_Kernel34_Valid_Out & channel20_Kernel34_Valid_Out & channel21_Kernel34_Valid_Out & channel22_Kernel34_Valid_Out & channel23_Kernel34_Valid_Out & channel24_Kernel34_Valid_Out & channel25_Kernel34_Valid_Out & channel26_Kernel34_Valid_Out & channel27_Kernel34_Valid_Out & channel28_Kernel34_Valid_Out & channel29_Kernel34_Valid_Out & channel30_Kernel34_Valid_Out & channel31_Kernel34_Valid_Out & channel32_Kernel34_Valid_Out & channel33_Kernel34_Valid_Out & channel34_Kernel34_Valid_Out & channel35_Kernel34_Valid_Out & channel36_Kernel34_Valid_Out & channel37_Kernel34_Valid_Out & channel38_Kernel34_Valid_Out & channel39_Kernel34_Valid_Out & channel40_Kernel34_Valid_Out & channel41_Kernel34_Valid_Out & channel42_Kernel34_Valid_Out & channel43_Kernel34_Valid_Out & channel44_Kernel34_Valid_Out & channel45_Kernel34_Valid_Out & channel46_Kernel34_Valid_Out & channel47_Kernel34_Valid_Out & channel48_Kernel34_Valid_Out & channel49_Kernel34_Valid_Out & channel50_Kernel34_Valid_Out & channel51_Kernel34_Valid_Out & channel52_Kernel34_Valid_Out & channel53_Kernel34_Valid_Out & channel54_Kernel34_Valid_Out & channel55_Kernel34_Valid_Out & channel56_Kernel34_Valid_Out & channel57_Kernel34_Valid_Out & channel58_Kernel34_Valid_Out & channel59_Kernel34_Valid_Out & channel60_Kernel34_Valid_Out & channel61_Kernel34_Valid_Out & channel62_Kernel34_Valid_Out & channel63_Kernel34_Valid_Out & channel64_Kernel34_Valid_Out;

	wire channel1_Kernel35_Valid_Out, channel2_Kernel35_Valid_Out, channel3_Kernel35_Valid_Out, channel4_Kernel35_Valid_Out, channel5_Kernel35_Valid_Out, channel6_Kernel35_Valid_Out, channel7_Kernel35_Valid_Out, channel8_Kernel35_Valid_Out, channel9_Kernel35_Valid_Out, channel10_Kernel35_Valid_Out, channel11_Kernel35_Valid_Out, channel12_Kernel35_Valid_Out, channel13_Kernel35_Valid_Out, channel14_Kernel35_Valid_Out, channel15_Kernel35_Valid_Out, channel16_Kernel35_Valid_Out, channel17_Kernel35_Valid_Out, channel18_Kernel35_Valid_Out, channel19_Kernel35_Valid_Out, channel20_Kernel35_Valid_Out, channel21_Kernel35_Valid_Out, channel22_Kernel35_Valid_Out, channel23_Kernel35_Valid_Out, channel24_Kernel35_Valid_Out, channel25_Kernel35_Valid_Out, channel26_Kernel35_Valid_Out, channel27_Kernel35_Valid_Out, channel28_Kernel35_Valid_Out, channel29_Kernel35_Valid_Out, channel30_Kernel35_Valid_Out, channel31_Kernel35_Valid_Out, channel32_Kernel35_Valid_Out, channel33_Kernel35_Valid_Out, channel34_Kernel35_Valid_Out, channel35_Kernel35_Valid_Out, channel36_Kernel35_Valid_Out, channel37_Kernel35_Valid_Out, channel38_Kernel35_Valid_Out, channel39_Kernel35_Valid_Out, channel40_Kernel35_Valid_Out, channel41_Kernel35_Valid_Out, channel42_Kernel35_Valid_Out, channel43_Kernel35_Valid_Out, channel44_Kernel35_Valid_Out, channel45_Kernel35_Valid_Out, channel46_Kernel35_Valid_Out, channel47_Kernel35_Valid_Out, channel48_Kernel35_Valid_Out, channel49_Kernel35_Valid_Out, channel50_Kernel35_Valid_Out, channel51_Kernel35_Valid_Out, channel52_Kernel35_Valid_Out, channel53_Kernel35_Valid_Out, channel54_Kernel35_Valid_Out, channel55_Kernel35_Valid_Out, channel56_Kernel35_Valid_Out, channel57_Kernel35_Valid_Out, channel58_Kernel35_Valid_Out, channel59_Kernel35_Valid_Out, channel60_Kernel35_Valid_Out, channel61_Kernel35_Valid_Out, channel62_Kernel35_Valid_Out, channel63_Kernel35_Valid_Out, channel64_Kernel35_Valid_Out;

	assign add_kernel35=channel1_Kernel35_Valid_Out & channel2_Kernel35_Valid_Out & channel3_Kernel35_Valid_Out & channel4_Kernel35_Valid_Out & channel5_Kernel35_Valid_Out & channel6_Kernel35_Valid_Out & channel7_Kernel35_Valid_Out & channel8_Kernel35_Valid_Out & channel9_Kernel35_Valid_Out & channel10_Kernel35_Valid_Out & channel11_Kernel35_Valid_Out & channel12_Kernel35_Valid_Out & channel13_Kernel35_Valid_Out & channel14_Kernel35_Valid_Out & channel15_Kernel35_Valid_Out & channel16_Kernel35_Valid_Out & channel17_Kernel35_Valid_Out & channel18_Kernel35_Valid_Out & channel19_Kernel35_Valid_Out & channel20_Kernel35_Valid_Out & channel21_Kernel35_Valid_Out & channel22_Kernel35_Valid_Out & channel23_Kernel35_Valid_Out & channel24_Kernel35_Valid_Out & channel25_Kernel35_Valid_Out & channel26_Kernel35_Valid_Out & channel27_Kernel35_Valid_Out & channel28_Kernel35_Valid_Out & channel29_Kernel35_Valid_Out & channel30_Kernel35_Valid_Out & channel31_Kernel35_Valid_Out & channel32_Kernel35_Valid_Out & channel33_Kernel35_Valid_Out & channel34_Kernel35_Valid_Out & channel35_Kernel35_Valid_Out & channel36_Kernel35_Valid_Out & channel37_Kernel35_Valid_Out & channel38_Kernel35_Valid_Out & channel39_Kernel35_Valid_Out & channel40_Kernel35_Valid_Out & channel41_Kernel35_Valid_Out & channel42_Kernel35_Valid_Out & channel43_Kernel35_Valid_Out & channel44_Kernel35_Valid_Out & channel45_Kernel35_Valid_Out & channel46_Kernel35_Valid_Out & channel47_Kernel35_Valid_Out & channel48_Kernel35_Valid_Out & channel49_Kernel35_Valid_Out & channel50_Kernel35_Valid_Out & channel51_Kernel35_Valid_Out & channel52_Kernel35_Valid_Out & channel53_Kernel35_Valid_Out & channel54_Kernel35_Valid_Out & channel55_Kernel35_Valid_Out & channel56_Kernel35_Valid_Out & channel57_Kernel35_Valid_Out & channel58_Kernel35_Valid_Out & channel59_Kernel35_Valid_Out & channel60_Kernel35_Valid_Out & channel61_Kernel35_Valid_Out & channel62_Kernel35_Valid_Out & channel63_Kernel35_Valid_Out & channel64_Kernel35_Valid_Out;

	wire channel1_Kernel36_Valid_Out, channel2_Kernel36_Valid_Out, channel3_Kernel36_Valid_Out, channel4_Kernel36_Valid_Out, channel5_Kernel36_Valid_Out, channel6_Kernel36_Valid_Out, channel7_Kernel36_Valid_Out, channel8_Kernel36_Valid_Out, channel9_Kernel36_Valid_Out, channel10_Kernel36_Valid_Out, channel11_Kernel36_Valid_Out, channel12_Kernel36_Valid_Out, channel13_Kernel36_Valid_Out, channel14_Kernel36_Valid_Out, channel15_Kernel36_Valid_Out, channel16_Kernel36_Valid_Out, channel17_Kernel36_Valid_Out, channel18_Kernel36_Valid_Out, channel19_Kernel36_Valid_Out, channel20_Kernel36_Valid_Out, channel21_Kernel36_Valid_Out, channel22_Kernel36_Valid_Out, channel23_Kernel36_Valid_Out, channel24_Kernel36_Valid_Out, channel25_Kernel36_Valid_Out, channel26_Kernel36_Valid_Out, channel27_Kernel36_Valid_Out, channel28_Kernel36_Valid_Out, channel29_Kernel36_Valid_Out, channel30_Kernel36_Valid_Out, channel31_Kernel36_Valid_Out, channel32_Kernel36_Valid_Out, channel33_Kernel36_Valid_Out, channel34_Kernel36_Valid_Out, channel35_Kernel36_Valid_Out, channel36_Kernel36_Valid_Out, channel37_Kernel36_Valid_Out, channel38_Kernel36_Valid_Out, channel39_Kernel36_Valid_Out, channel40_Kernel36_Valid_Out, channel41_Kernel36_Valid_Out, channel42_Kernel36_Valid_Out, channel43_Kernel36_Valid_Out, channel44_Kernel36_Valid_Out, channel45_Kernel36_Valid_Out, channel46_Kernel36_Valid_Out, channel47_Kernel36_Valid_Out, channel48_Kernel36_Valid_Out, channel49_Kernel36_Valid_Out, channel50_Kernel36_Valid_Out, channel51_Kernel36_Valid_Out, channel52_Kernel36_Valid_Out, channel53_Kernel36_Valid_Out, channel54_Kernel36_Valid_Out, channel55_Kernel36_Valid_Out, channel56_Kernel36_Valid_Out, channel57_Kernel36_Valid_Out, channel58_Kernel36_Valid_Out, channel59_Kernel36_Valid_Out, channel60_Kernel36_Valid_Out, channel61_Kernel36_Valid_Out, channel62_Kernel36_Valid_Out, channel63_Kernel36_Valid_Out, channel64_Kernel36_Valid_Out;

	assign add_kernel36=channel1_Kernel36_Valid_Out & channel2_Kernel36_Valid_Out & channel3_Kernel36_Valid_Out & channel4_Kernel36_Valid_Out & channel5_Kernel36_Valid_Out & channel6_Kernel36_Valid_Out & channel7_Kernel36_Valid_Out & channel8_Kernel36_Valid_Out & channel9_Kernel36_Valid_Out & channel10_Kernel36_Valid_Out & channel11_Kernel36_Valid_Out & channel12_Kernel36_Valid_Out & channel13_Kernel36_Valid_Out & channel14_Kernel36_Valid_Out & channel15_Kernel36_Valid_Out & channel16_Kernel36_Valid_Out & channel17_Kernel36_Valid_Out & channel18_Kernel36_Valid_Out & channel19_Kernel36_Valid_Out & channel20_Kernel36_Valid_Out & channel21_Kernel36_Valid_Out & channel22_Kernel36_Valid_Out & channel23_Kernel36_Valid_Out & channel24_Kernel36_Valid_Out & channel25_Kernel36_Valid_Out & channel26_Kernel36_Valid_Out & channel27_Kernel36_Valid_Out & channel28_Kernel36_Valid_Out & channel29_Kernel36_Valid_Out & channel30_Kernel36_Valid_Out & channel31_Kernel36_Valid_Out & channel32_Kernel36_Valid_Out & channel33_Kernel36_Valid_Out & channel34_Kernel36_Valid_Out & channel35_Kernel36_Valid_Out & channel36_Kernel36_Valid_Out & channel37_Kernel36_Valid_Out & channel38_Kernel36_Valid_Out & channel39_Kernel36_Valid_Out & channel40_Kernel36_Valid_Out & channel41_Kernel36_Valid_Out & channel42_Kernel36_Valid_Out & channel43_Kernel36_Valid_Out & channel44_Kernel36_Valid_Out & channel45_Kernel36_Valid_Out & channel46_Kernel36_Valid_Out & channel47_Kernel36_Valid_Out & channel48_Kernel36_Valid_Out & channel49_Kernel36_Valid_Out & channel50_Kernel36_Valid_Out & channel51_Kernel36_Valid_Out & channel52_Kernel36_Valid_Out & channel53_Kernel36_Valid_Out & channel54_Kernel36_Valid_Out & channel55_Kernel36_Valid_Out & channel56_Kernel36_Valid_Out & channel57_Kernel36_Valid_Out & channel58_Kernel36_Valid_Out & channel59_Kernel36_Valid_Out & channel60_Kernel36_Valid_Out & channel61_Kernel36_Valid_Out & channel62_Kernel36_Valid_Out & channel63_Kernel36_Valid_Out & channel64_Kernel36_Valid_Out;

	wire channel1_Kernel37_Valid_Out, channel2_Kernel37_Valid_Out, channel3_Kernel37_Valid_Out, channel4_Kernel37_Valid_Out, channel5_Kernel37_Valid_Out, channel6_Kernel37_Valid_Out, channel7_Kernel37_Valid_Out, channel8_Kernel37_Valid_Out, channel9_Kernel37_Valid_Out, channel10_Kernel37_Valid_Out, channel11_Kernel37_Valid_Out, channel12_Kernel37_Valid_Out, channel13_Kernel37_Valid_Out, channel14_Kernel37_Valid_Out, channel15_Kernel37_Valid_Out, channel16_Kernel37_Valid_Out, channel17_Kernel37_Valid_Out, channel18_Kernel37_Valid_Out, channel19_Kernel37_Valid_Out, channel20_Kernel37_Valid_Out, channel21_Kernel37_Valid_Out, channel22_Kernel37_Valid_Out, channel23_Kernel37_Valid_Out, channel24_Kernel37_Valid_Out, channel25_Kernel37_Valid_Out, channel26_Kernel37_Valid_Out, channel27_Kernel37_Valid_Out, channel28_Kernel37_Valid_Out, channel29_Kernel37_Valid_Out, channel30_Kernel37_Valid_Out, channel31_Kernel37_Valid_Out, channel32_Kernel37_Valid_Out, channel33_Kernel37_Valid_Out, channel34_Kernel37_Valid_Out, channel35_Kernel37_Valid_Out, channel36_Kernel37_Valid_Out, channel37_Kernel37_Valid_Out, channel38_Kernel37_Valid_Out, channel39_Kernel37_Valid_Out, channel40_Kernel37_Valid_Out, channel41_Kernel37_Valid_Out, channel42_Kernel37_Valid_Out, channel43_Kernel37_Valid_Out, channel44_Kernel37_Valid_Out, channel45_Kernel37_Valid_Out, channel46_Kernel37_Valid_Out, channel47_Kernel37_Valid_Out, channel48_Kernel37_Valid_Out, channel49_Kernel37_Valid_Out, channel50_Kernel37_Valid_Out, channel51_Kernel37_Valid_Out, channel52_Kernel37_Valid_Out, channel53_Kernel37_Valid_Out, channel54_Kernel37_Valid_Out, channel55_Kernel37_Valid_Out, channel56_Kernel37_Valid_Out, channel57_Kernel37_Valid_Out, channel58_Kernel37_Valid_Out, channel59_Kernel37_Valid_Out, channel60_Kernel37_Valid_Out, channel61_Kernel37_Valid_Out, channel62_Kernel37_Valid_Out, channel63_Kernel37_Valid_Out, channel64_Kernel37_Valid_Out;

	assign add_kernel37=channel1_Kernel37_Valid_Out & channel2_Kernel37_Valid_Out & channel3_Kernel37_Valid_Out & channel4_Kernel37_Valid_Out & channel5_Kernel37_Valid_Out & channel6_Kernel37_Valid_Out & channel7_Kernel37_Valid_Out & channel8_Kernel37_Valid_Out & channel9_Kernel37_Valid_Out & channel10_Kernel37_Valid_Out & channel11_Kernel37_Valid_Out & channel12_Kernel37_Valid_Out & channel13_Kernel37_Valid_Out & channel14_Kernel37_Valid_Out & channel15_Kernel37_Valid_Out & channel16_Kernel37_Valid_Out & channel17_Kernel37_Valid_Out & channel18_Kernel37_Valid_Out & channel19_Kernel37_Valid_Out & channel20_Kernel37_Valid_Out & channel21_Kernel37_Valid_Out & channel22_Kernel37_Valid_Out & channel23_Kernel37_Valid_Out & channel24_Kernel37_Valid_Out & channel25_Kernel37_Valid_Out & channel26_Kernel37_Valid_Out & channel27_Kernel37_Valid_Out & channel28_Kernel37_Valid_Out & channel29_Kernel37_Valid_Out & channel30_Kernel37_Valid_Out & channel31_Kernel37_Valid_Out & channel32_Kernel37_Valid_Out & channel33_Kernel37_Valid_Out & channel34_Kernel37_Valid_Out & channel35_Kernel37_Valid_Out & channel36_Kernel37_Valid_Out & channel37_Kernel37_Valid_Out & channel38_Kernel37_Valid_Out & channel39_Kernel37_Valid_Out & channel40_Kernel37_Valid_Out & channel41_Kernel37_Valid_Out & channel42_Kernel37_Valid_Out & channel43_Kernel37_Valid_Out & channel44_Kernel37_Valid_Out & channel45_Kernel37_Valid_Out & channel46_Kernel37_Valid_Out & channel47_Kernel37_Valid_Out & channel48_Kernel37_Valid_Out & channel49_Kernel37_Valid_Out & channel50_Kernel37_Valid_Out & channel51_Kernel37_Valid_Out & channel52_Kernel37_Valid_Out & channel53_Kernel37_Valid_Out & channel54_Kernel37_Valid_Out & channel55_Kernel37_Valid_Out & channel56_Kernel37_Valid_Out & channel57_Kernel37_Valid_Out & channel58_Kernel37_Valid_Out & channel59_Kernel37_Valid_Out & channel60_Kernel37_Valid_Out & channel61_Kernel37_Valid_Out & channel62_Kernel37_Valid_Out & channel63_Kernel37_Valid_Out & channel64_Kernel37_Valid_Out;

	wire channel1_Kernel38_Valid_Out, channel2_Kernel38_Valid_Out, channel3_Kernel38_Valid_Out, channel4_Kernel38_Valid_Out, channel5_Kernel38_Valid_Out, channel6_Kernel38_Valid_Out, channel7_Kernel38_Valid_Out, channel8_Kernel38_Valid_Out, channel9_Kernel38_Valid_Out, channel10_Kernel38_Valid_Out, channel11_Kernel38_Valid_Out, channel12_Kernel38_Valid_Out, channel13_Kernel38_Valid_Out, channel14_Kernel38_Valid_Out, channel15_Kernel38_Valid_Out, channel16_Kernel38_Valid_Out, channel17_Kernel38_Valid_Out, channel18_Kernel38_Valid_Out, channel19_Kernel38_Valid_Out, channel20_Kernel38_Valid_Out, channel21_Kernel38_Valid_Out, channel22_Kernel38_Valid_Out, channel23_Kernel38_Valid_Out, channel24_Kernel38_Valid_Out, channel25_Kernel38_Valid_Out, channel26_Kernel38_Valid_Out, channel27_Kernel38_Valid_Out, channel28_Kernel38_Valid_Out, channel29_Kernel38_Valid_Out, channel30_Kernel38_Valid_Out, channel31_Kernel38_Valid_Out, channel32_Kernel38_Valid_Out, channel33_Kernel38_Valid_Out, channel34_Kernel38_Valid_Out, channel35_Kernel38_Valid_Out, channel36_Kernel38_Valid_Out, channel37_Kernel38_Valid_Out, channel38_Kernel38_Valid_Out, channel39_Kernel38_Valid_Out, channel40_Kernel38_Valid_Out, channel41_Kernel38_Valid_Out, channel42_Kernel38_Valid_Out, channel43_Kernel38_Valid_Out, channel44_Kernel38_Valid_Out, channel45_Kernel38_Valid_Out, channel46_Kernel38_Valid_Out, channel47_Kernel38_Valid_Out, channel48_Kernel38_Valid_Out, channel49_Kernel38_Valid_Out, channel50_Kernel38_Valid_Out, channel51_Kernel38_Valid_Out, channel52_Kernel38_Valid_Out, channel53_Kernel38_Valid_Out, channel54_Kernel38_Valid_Out, channel55_Kernel38_Valid_Out, channel56_Kernel38_Valid_Out, channel57_Kernel38_Valid_Out, channel58_Kernel38_Valid_Out, channel59_Kernel38_Valid_Out, channel60_Kernel38_Valid_Out, channel61_Kernel38_Valid_Out, channel62_Kernel38_Valid_Out, channel63_Kernel38_Valid_Out, channel64_Kernel38_Valid_Out;

	assign add_kernel38=channel1_Kernel38_Valid_Out & channel2_Kernel38_Valid_Out & channel3_Kernel38_Valid_Out & channel4_Kernel38_Valid_Out & channel5_Kernel38_Valid_Out & channel6_Kernel38_Valid_Out & channel7_Kernel38_Valid_Out & channel8_Kernel38_Valid_Out & channel9_Kernel38_Valid_Out & channel10_Kernel38_Valid_Out & channel11_Kernel38_Valid_Out & channel12_Kernel38_Valid_Out & channel13_Kernel38_Valid_Out & channel14_Kernel38_Valid_Out & channel15_Kernel38_Valid_Out & channel16_Kernel38_Valid_Out & channel17_Kernel38_Valid_Out & channel18_Kernel38_Valid_Out & channel19_Kernel38_Valid_Out & channel20_Kernel38_Valid_Out & channel21_Kernel38_Valid_Out & channel22_Kernel38_Valid_Out & channel23_Kernel38_Valid_Out & channel24_Kernel38_Valid_Out & channel25_Kernel38_Valid_Out & channel26_Kernel38_Valid_Out & channel27_Kernel38_Valid_Out & channel28_Kernel38_Valid_Out & channel29_Kernel38_Valid_Out & channel30_Kernel38_Valid_Out & channel31_Kernel38_Valid_Out & channel32_Kernel38_Valid_Out & channel33_Kernel38_Valid_Out & channel34_Kernel38_Valid_Out & channel35_Kernel38_Valid_Out & channel36_Kernel38_Valid_Out & channel37_Kernel38_Valid_Out & channel38_Kernel38_Valid_Out & channel39_Kernel38_Valid_Out & channel40_Kernel38_Valid_Out & channel41_Kernel38_Valid_Out & channel42_Kernel38_Valid_Out & channel43_Kernel38_Valid_Out & channel44_Kernel38_Valid_Out & channel45_Kernel38_Valid_Out & channel46_Kernel38_Valid_Out & channel47_Kernel38_Valid_Out & channel48_Kernel38_Valid_Out & channel49_Kernel38_Valid_Out & channel50_Kernel38_Valid_Out & channel51_Kernel38_Valid_Out & channel52_Kernel38_Valid_Out & channel53_Kernel38_Valid_Out & channel54_Kernel38_Valid_Out & channel55_Kernel38_Valid_Out & channel56_Kernel38_Valid_Out & channel57_Kernel38_Valid_Out & channel58_Kernel38_Valid_Out & channel59_Kernel38_Valid_Out & channel60_Kernel38_Valid_Out & channel61_Kernel38_Valid_Out & channel62_Kernel38_Valid_Out & channel63_Kernel38_Valid_Out & channel64_Kernel38_Valid_Out;

	wire channel1_Kernel39_Valid_Out, channel2_Kernel39_Valid_Out, channel3_Kernel39_Valid_Out, channel4_Kernel39_Valid_Out, channel5_Kernel39_Valid_Out, channel6_Kernel39_Valid_Out, channel7_Kernel39_Valid_Out, channel8_Kernel39_Valid_Out, channel9_Kernel39_Valid_Out, channel10_Kernel39_Valid_Out, channel11_Kernel39_Valid_Out, channel12_Kernel39_Valid_Out, channel13_Kernel39_Valid_Out, channel14_Kernel39_Valid_Out, channel15_Kernel39_Valid_Out, channel16_Kernel39_Valid_Out, channel17_Kernel39_Valid_Out, channel18_Kernel39_Valid_Out, channel19_Kernel39_Valid_Out, channel20_Kernel39_Valid_Out, channel21_Kernel39_Valid_Out, channel22_Kernel39_Valid_Out, channel23_Kernel39_Valid_Out, channel24_Kernel39_Valid_Out, channel25_Kernel39_Valid_Out, channel26_Kernel39_Valid_Out, channel27_Kernel39_Valid_Out, channel28_Kernel39_Valid_Out, channel29_Kernel39_Valid_Out, channel30_Kernel39_Valid_Out, channel31_Kernel39_Valid_Out, channel32_Kernel39_Valid_Out, channel33_Kernel39_Valid_Out, channel34_Kernel39_Valid_Out, channel35_Kernel39_Valid_Out, channel36_Kernel39_Valid_Out, channel37_Kernel39_Valid_Out, channel38_Kernel39_Valid_Out, channel39_Kernel39_Valid_Out, channel40_Kernel39_Valid_Out, channel41_Kernel39_Valid_Out, channel42_Kernel39_Valid_Out, channel43_Kernel39_Valid_Out, channel44_Kernel39_Valid_Out, channel45_Kernel39_Valid_Out, channel46_Kernel39_Valid_Out, channel47_Kernel39_Valid_Out, channel48_Kernel39_Valid_Out, channel49_Kernel39_Valid_Out, channel50_Kernel39_Valid_Out, channel51_Kernel39_Valid_Out, channel52_Kernel39_Valid_Out, channel53_Kernel39_Valid_Out, channel54_Kernel39_Valid_Out, channel55_Kernel39_Valid_Out, channel56_Kernel39_Valid_Out, channel57_Kernel39_Valid_Out, channel58_Kernel39_Valid_Out, channel59_Kernel39_Valid_Out, channel60_Kernel39_Valid_Out, channel61_Kernel39_Valid_Out, channel62_Kernel39_Valid_Out, channel63_Kernel39_Valid_Out, channel64_Kernel39_Valid_Out;

	assign add_kernel39=channel1_Kernel39_Valid_Out & channel2_Kernel39_Valid_Out & channel3_Kernel39_Valid_Out & channel4_Kernel39_Valid_Out & channel5_Kernel39_Valid_Out & channel6_Kernel39_Valid_Out & channel7_Kernel39_Valid_Out & channel8_Kernel39_Valid_Out & channel9_Kernel39_Valid_Out & channel10_Kernel39_Valid_Out & channel11_Kernel39_Valid_Out & channel12_Kernel39_Valid_Out & channel13_Kernel39_Valid_Out & channel14_Kernel39_Valid_Out & channel15_Kernel39_Valid_Out & channel16_Kernel39_Valid_Out & channel17_Kernel39_Valid_Out & channel18_Kernel39_Valid_Out & channel19_Kernel39_Valid_Out & channel20_Kernel39_Valid_Out & channel21_Kernel39_Valid_Out & channel22_Kernel39_Valid_Out & channel23_Kernel39_Valid_Out & channel24_Kernel39_Valid_Out & channel25_Kernel39_Valid_Out & channel26_Kernel39_Valid_Out & channel27_Kernel39_Valid_Out & channel28_Kernel39_Valid_Out & channel29_Kernel39_Valid_Out & channel30_Kernel39_Valid_Out & channel31_Kernel39_Valid_Out & channel32_Kernel39_Valid_Out & channel33_Kernel39_Valid_Out & channel34_Kernel39_Valid_Out & channel35_Kernel39_Valid_Out & channel36_Kernel39_Valid_Out & channel37_Kernel39_Valid_Out & channel38_Kernel39_Valid_Out & channel39_Kernel39_Valid_Out & channel40_Kernel39_Valid_Out & channel41_Kernel39_Valid_Out & channel42_Kernel39_Valid_Out & channel43_Kernel39_Valid_Out & channel44_Kernel39_Valid_Out & channel45_Kernel39_Valid_Out & channel46_Kernel39_Valid_Out & channel47_Kernel39_Valid_Out & channel48_Kernel39_Valid_Out & channel49_Kernel39_Valid_Out & channel50_Kernel39_Valid_Out & channel51_Kernel39_Valid_Out & channel52_Kernel39_Valid_Out & channel53_Kernel39_Valid_Out & channel54_Kernel39_Valid_Out & channel55_Kernel39_Valid_Out & channel56_Kernel39_Valid_Out & channel57_Kernel39_Valid_Out & channel58_Kernel39_Valid_Out & channel59_Kernel39_Valid_Out & channel60_Kernel39_Valid_Out & channel61_Kernel39_Valid_Out & channel62_Kernel39_Valid_Out & channel63_Kernel39_Valid_Out & channel64_Kernel39_Valid_Out;

	wire channel1_Kernel40_Valid_Out, channel2_Kernel40_Valid_Out, channel3_Kernel40_Valid_Out, channel4_Kernel40_Valid_Out, channel5_Kernel40_Valid_Out, channel6_Kernel40_Valid_Out, channel7_Kernel40_Valid_Out, channel8_Kernel40_Valid_Out, channel9_Kernel40_Valid_Out, channel10_Kernel40_Valid_Out, channel11_Kernel40_Valid_Out, channel12_Kernel40_Valid_Out, channel13_Kernel40_Valid_Out, channel14_Kernel40_Valid_Out, channel15_Kernel40_Valid_Out, channel16_Kernel40_Valid_Out, channel17_Kernel40_Valid_Out, channel18_Kernel40_Valid_Out, channel19_Kernel40_Valid_Out, channel20_Kernel40_Valid_Out, channel21_Kernel40_Valid_Out, channel22_Kernel40_Valid_Out, channel23_Kernel40_Valid_Out, channel24_Kernel40_Valid_Out, channel25_Kernel40_Valid_Out, channel26_Kernel40_Valid_Out, channel27_Kernel40_Valid_Out, channel28_Kernel40_Valid_Out, channel29_Kernel40_Valid_Out, channel30_Kernel40_Valid_Out, channel31_Kernel40_Valid_Out, channel32_Kernel40_Valid_Out, channel33_Kernel40_Valid_Out, channel34_Kernel40_Valid_Out, channel35_Kernel40_Valid_Out, channel36_Kernel40_Valid_Out, channel37_Kernel40_Valid_Out, channel38_Kernel40_Valid_Out, channel39_Kernel40_Valid_Out, channel40_Kernel40_Valid_Out, channel41_Kernel40_Valid_Out, channel42_Kernel40_Valid_Out, channel43_Kernel40_Valid_Out, channel44_Kernel40_Valid_Out, channel45_Kernel40_Valid_Out, channel46_Kernel40_Valid_Out, channel47_Kernel40_Valid_Out, channel48_Kernel40_Valid_Out, channel49_Kernel40_Valid_Out, channel50_Kernel40_Valid_Out, channel51_Kernel40_Valid_Out, channel52_Kernel40_Valid_Out, channel53_Kernel40_Valid_Out, channel54_Kernel40_Valid_Out, channel55_Kernel40_Valid_Out, channel56_Kernel40_Valid_Out, channel57_Kernel40_Valid_Out, channel58_Kernel40_Valid_Out, channel59_Kernel40_Valid_Out, channel60_Kernel40_Valid_Out, channel61_Kernel40_Valid_Out, channel62_Kernel40_Valid_Out, channel63_Kernel40_Valid_Out, channel64_Kernel40_Valid_Out;

	assign add_kernel40=channel1_Kernel40_Valid_Out & channel2_Kernel40_Valid_Out & channel3_Kernel40_Valid_Out & channel4_Kernel40_Valid_Out & channel5_Kernel40_Valid_Out & channel6_Kernel40_Valid_Out & channel7_Kernel40_Valid_Out & channel8_Kernel40_Valid_Out & channel9_Kernel40_Valid_Out & channel10_Kernel40_Valid_Out & channel11_Kernel40_Valid_Out & channel12_Kernel40_Valid_Out & channel13_Kernel40_Valid_Out & channel14_Kernel40_Valid_Out & channel15_Kernel40_Valid_Out & channel16_Kernel40_Valid_Out & channel17_Kernel40_Valid_Out & channel18_Kernel40_Valid_Out & channel19_Kernel40_Valid_Out & channel20_Kernel40_Valid_Out & channel21_Kernel40_Valid_Out & channel22_Kernel40_Valid_Out & channel23_Kernel40_Valid_Out & channel24_Kernel40_Valid_Out & channel25_Kernel40_Valid_Out & channel26_Kernel40_Valid_Out & channel27_Kernel40_Valid_Out & channel28_Kernel40_Valid_Out & channel29_Kernel40_Valid_Out & channel30_Kernel40_Valid_Out & channel31_Kernel40_Valid_Out & channel32_Kernel40_Valid_Out & channel33_Kernel40_Valid_Out & channel34_Kernel40_Valid_Out & channel35_Kernel40_Valid_Out & channel36_Kernel40_Valid_Out & channel37_Kernel40_Valid_Out & channel38_Kernel40_Valid_Out & channel39_Kernel40_Valid_Out & channel40_Kernel40_Valid_Out & channel41_Kernel40_Valid_Out & channel42_Kernel40_Valid_Out & channel43_Kernel40_Valid_Out & channel44_Kernel40_Valid_Out & channel45_Kernel40_Valid_Out & channel46_Kernel40_Valid_Out & channel47_Kernel40_Valid_Out & channel48_Kernel40_Valid_Out & channel49_Kernel40_Valid_Out & channel50_Kernel40_Valid_Out & channel51_Kernel40_Valid_Out & channel52_Kernel40_Valid_Out & channel53_Kernel40_Valid_Out & channel54_Kernel40_Valid_Out & channel55_Kernel40_Valid_Out & channel56_Kernel40_Valid_Out & channel57_Kernel40_Valid_Out & channel58_Kernel40_Valid_Out & channel59_Kernel40_Valid_Out & channel60_Kernel40_Valid_Out & channel61_Kernel40_Valid_Out & channel62_Kernel40_Valid_Out & channel63_Kernel40_Valid_Out & channel64_Kernel40_Valid_Out;

	wire channel1_Kernel41_Valid_Out, channel2_Kernel41_Valid_Out, channel3_Kernel41_Valid_Out, channel4_Kernel41_Valid_Out, channel5_Kernel41_Valid_Out, channel6_Kernel41_Valid_Out, channel7_Kernel41_Valid_Out, channel8_Kernel41_Valid_Out, channel9_Kernel41_Valid_Out, channel10_Kernel41_Valid_Out, channel11_Kernel41_Valid_Out, channel12_Kernel41_Valid_Out, channel13_Kernel41_Valid_Out, channel14_Kernel41_Valid_Out, channel15_Kernel41_Valid_Out, channel16_Kernel41_Valid_Out, channel17_Kernel41_Valid_Out, channel18_Kernel41_Valid_Out, channel19_Kernel41_Valid_Out, channel20_Kernel41_Valid_Out, channel21_Kernel41_Valid_Out, channel22_Kernel41_Valid_Out, channel23_Kernel41_Valid_Out, channel24_Kernel41_Valid_Out, channel25_Kernel41_Valid_Out, channel26_Kernel41_Valid_Out, channel27_Kernel41_Valid_Out, channel28_Kernel41_Valid_Out, channel29_Kernel41_Valid_Out, channel30_Kernel41_Valid_Out, channel31_Kernel41_Valid_Out, channel32_Kernel41_Valid_Out, channel33_Kernel41_Valid_Out, channel34_Kernel41_Valid_Out, channel35_Kernel41_Valid_Out, channel36_Kernel41_Valid_Out, channel37_Kernel41_Valid_Out, channel38_Kernel41_Valid_Out, channel39_Kernel41_Valid_Out, channel40_Kernel41_Valid_Out, channel41_Kernel41_Valid_Out, channel42_Kernel41_Valid_Out, channel43_Kernel41_Valid_Out, channel44_Kernel41_Valid_Out, channel45_Kernel41_Valid_Out, channel46_Kernel41_Valid_Out, channel47_Kernel41_Valid_Out, channel48_Kernel41_Valid_Out, channel49_Kernel41_Valid_Out, channel50_Kernel41_Valid_Out, channel51_Kernel41_Valid_Out, channel52_Kernel41_Valid_Out, channel53_Kernel41_Valid_Out, channel54_Kernel41_Valid_Out, channel55_Kernel41_Valid_Out, channel56_Kernel41_Valid_Out, channel57_Kernel41_Valid_Out, channel58_Kernel41_Valid_Out, channel59_Kernel41_Valid_Out, channel60_Kernel41_Valid_Out, channel61_Kernel41_Valid_Out, channel62_Kernel41_Valid_Out, channel63_Kernel41_Valid_Out, channel64_Kernel41_Valid_Out;

	assign add_kernel41=channel1_Kernel41_Valid_Out & channel2_Kernel41_Valid_Out & channel3_Kernel41_Valid_Out & channel4_Kernel41_Valid_Out & channel5_Kernel41_Valid_Out & channel6_Kernel41_Valid_Out & channel7_Kernel41_Valid_Out & channel8_Kernel41_Valid_Out & channel9_Kernel41_Valid_Out & channel10_Kernel41_Valid_Out & channel11_Kernel41_Valid_Out & channel12_Kernel41_Valid_Out & channel13_Kernel41_Valid_Out & channel14_Kernel41_Valid_Out & channel15_Kernel41_Valid_Out & channel16_Kernel41_Valid_Out & channel17_Kernel41_Valid_Out & channel18_Kernel41_Valid_Out & channel19_Kernel41_Valid_Out & channel20_Kernel41_Valid_Out & channel21_Kernel41_Valid_Out & channel22_Kernel41_Valid_Out & channel23_Kernel41_Valid_Out & channel24_Kernel41_Valid_Out & channel25_Kernel41_Valid_Out & channel26_Kernel41_Valid_Out & channel27_Kernel41_Valid_Out & channel28_Kernel41_Valid_Out & channel29_Kernel41_Valid_Out & channel30_Kernel41_Valid_Out & channel31_Kernel41_Valid_Out & channel32_Kernel41_Valid_Out & channel33_Kernel41_Valid_Out & channel34_Kernel41_Valid_Out & channel35_Kernel41_Valid_Out & channel36_Kernel41_Valid_Out & channel37_Kernel41_Valid_Out & channel38_Kernel41_Valid_Out & channel39_Kernel41_Valid_Out & channel40_Kernel41_Valid_Out & channel41_Kernel41_Valid_Out & channel42_Kernel41_Valid_Out & channel43_Kernel41_Valid_Out & channel44_Kernel41_Valid_Out & channel45_Kernel41_Valid_Out & channel46_Kernel41_Valid_Out & channel47_Kernel41_Valid_Out & channel48_Kernel41_Valid_Out & channel49_Kernel41_Valid_Out & channel50_Kernel41_Valid_Out & channel51_Kernel41_Valid_Out & channel52_Kernel41_Valid_Out & channel53_Kernel41_Valid_Out & channel54_Kernel41_Valid_Out & channel55_Kernel41_Valid_Out & channel56_Kernel41_Valid_Out & channel57_Kernel41_Valid_Out & channel58_Kernel41_Valid_Out & channel59_Kernel41_Valid_Out & channel60_Kernel41_Valid_Out & channel61_Kernel41_Valid_Out & channel62_Kernel41_Valid_Out & channel63_Kernel41_Valid_Out & channel64_Kernel41_Valid_Out;

	wire channel1_Kernel42_Valid_Out, channel2_Kernel42_Valid_Out, channel3_Kernel42_Valid_Out, channel4_Kernel42_Valid_Out, channel5_Kernel42_Valid_Out, channel6_Kernel42_Valid_Out, channel7_Kernel42_Valid_Out, channel8_Kernel42_Valid_Out, channel9_Kernel42_Valid_Out, channel10_Kernel42_Valid_Out, channel11_Kernel42_Valid_Out, channel12_Kernel42_Valid_Out, channel13_Kernel42_Valid_Out, channel14_Kernel42_Valid_Out, channel15_Kernel42_Valid_Out, channel16_Kernel42_Valid_Out, channel17_Kernel42_Valid_Out, channel18_Kernel42_Valid_Out, channel19_Kernel42_Valid_Out, channel20_Kernel42_Valid_Out, channel21_Kernel42_Valid_Out, channel22_Kernel42_Valid_Out, channel23_Kernel42_Valid_Out, channel24_Kernel42_Valid_Out, channel25_Kernel42_Valid_Out, channel26_Kernel42_Valid_Out, channel27_Kernel42_Valid_Out, channel28_Kernel42_Valid_Out, channel29_Kernel42_Valid_Out, channel30_Kernel42_Valid_Out, channel31_Kernel42_Valid_Out, channel32_Kernel42_Valid_Out, channel33_Kernel42_Valid_Out, channel34_Kernel42_Valid_Out, channel35_Kernel42_Valid_Out, channel36_Kernel42_Valid_Out, channel37_Kernel42_Valid_Out, channel38_Kernel42_Valid_Out, channel39_Kernel42_Valid_Out, channel40_Kernel42_Valid_Out, channel41_Kernel42_Valid_Out, channel42_Kernel42_Valid_Out, channel43_Kernel42_Valid_Out, channel44_Kernel42_Valid_Out, channel45_Kernel42_Valid_Out, channel46_Kernel42_Valid_Out, channel47_Kernel42_Valid_Out, channel48_Kernel42_Valid_Out, channel49_Kernel42_Valid_Out, channel50_Kernel42_Valid_Out, channel51_Kernel42_Valid_Out, channel52_Kernel42_Valid_Out, channel53_Kernel42_Valid_Out, channel54_Kernel42_Valid_Out, channel55_Kernel42_Valid_Out, channel56_Kernel42_Valid_Out, channel57_Kernel42_Valid_Out, channel58_Kernel42_Valid_Out, channel59_Kernel42_Valid_Out, channel60_Kernel42_Valid_Out, channel61_Kernel42_Valid_Out, channel62_Kernel42_Valid_Out, channel63_Kernel42_Valid_Out, channel64_Kernel42_Valid_Out;

	assign add_kernel42=channel1_Kernel42_Valid_Out & channel2_Kernel42_Valid_Out & channel3_Kernel42_Valid_Out & channel4_Kernel42_Valid_Out & channel5_Kernel42_Valid_Out & channel6_Kernel42_Valid_Out & channel7_Kernel42_Valid_Out & channel8_Kernel42_Valid_Out & channel9_Kernel42_Valid_Out & channel10_Kernel42_Valid_Out & channel11_Kernel42_Valid_Out & channel12_Kernel42_Valid_Out & channel13_Kernel42_Valid_Out & channel14_Kernel42_Valid_Out & channel15_Kernel42_Valid_Out & channel16_Kernel42_Valid_Out & channel17_Kernel42_Valid_Out & channel18_Kernel42_Valid_Out & channel19_Kernel42_Valid_Out & channel20_Kernel42_Valid_Out & channel21_Kernel42_Valid_Out & channel22_Kernel42_Valid_Out & channel23_Kernel42_Valid_Out & channel24_Kernel42_Valid_Out & channel25_Kernel42_Valid_Out & channel26_Kernel42_Valid_Out & channel27_Kernel42_Valid_Out & channel28_Kernel42_Valid_Out & channel29_Kernel42_Valid_Out & channel30_Kernel42_Valid_Out & channel31_Kernel42_Valid_Out & channel32_Kernel42_Valid_Out & channel33_Kernel42_Valid_Out & channel34_Kernel42_Valid_Out & channel35_Kernel42_Valid_Out & channel36_Kernel42_Valid_Out & channel37_Kernel42_Valid_Out & channel38_Kernel42_Valid_Out & channel39_Kernel42_Valid_Out & channel40_Kernel42_Valid_Out & channel41_Kernel42_Valid_Out & channel42_Kernel42_Valid_Out & channel43_Kernel42_Valid_Out & channel44_Kernel42_Valid_Out & channel45_Kernel42_Valid_Out & channel46_Kernel42_Valid_Out & channel47_Kernel42_Valid_Out & channel48_Kernel42_Valid_Out & channel49_Kernel42_Valid_Out & channel50_Kernel42_Valid_Out & channel51_Kernel42_Valid_Out & channel52_Kernel42_Valid_Out & channel53_Kernel42_Valid_Out & channel54_Kernel42_Valid_Out & channel55_Kernel42_Valid_Out & channel56_Kernel42_Valid_Out & channel57_Kernel42_Valid_Out & channel58_Kernel42_Valid_Out & channel59_Kernel42_Valid_Out & channel60_Kernel42_Valid_Out & channel61_Kernel42_Valid_Out & channel62_Kernel42_Valid_Out & channel63_Kernel42_Valid_Out & channel64_Kernel42_Valid_Out;

	wire channel1_Kernel43_Valid_Out, channel2_Kernel43_Valid_Out, channel3_Kernel43_Valid_Out, channel4_Kernel43_Valid_Out, channel5_Kernel43_Valid_Out, channel6_Kernel43_Valid_Out, channel7_Kernel43_Valid_Out, channel8_Kernel43_Valid_Out, channel9_Kernel43_Valid_Out, channel10_Kernel43_Valid_Out, channel11_Kernel43_Valid_Out, channel12_Kernel43_Valid_Out, channel13_Kernel43_Valid_Out, channel14_Kernel43_Valid_Out, channel15_Kernel43_Valid_Out, channel16_Kernel43_Valid_Out, channel17_Kernel43_Valid_Out, channel18_Kernel43_Valid_Out, channel19_Kernel43_Valid_Out, channel20_Kernel43_Valid_Out, channel21_Kernel43_Valid_Out, channel22_Kernel43_Valid_Out, channel23_Kernel43_Valid_Out, channel24_Kernel43_Valid_Out, channel25_Kernel43_Valid_Out, channel26_Kernel43_Valid_Out, channel27_Kernel43_Valid_Out, channel28_Kernel43_Valid_Out, channel29_Kernel43_Valid_Out, channel30_Kernel43_Valid_Out, channel31_Kernel43_Valid_Out, channel32_Kernel43_Valid_Out, channel33_Kernel43_Valid_Out, channel34_Kernel43_Valid_Out, channel35_Kernel43_Valid_Out, channel36_Kernel43_Valid_Out, channel37_Kernel43_Valid_Out, channel38_Kernel43_Valid_Out, channel39_Kernel43_Valid_Out, channel40_Kernel43_Valid_Out, channel41_Kernel43_Valid_Out, channel42_Kernel43_Valid_Out, channel43_Kernel43_Valid_Out, channel44_Kernel43_Valid_Out, channel45_Kernel43_Valid_Out, channel46_Kernel43_Valid_Out, channel47_Kernel43_Valid_Out, channel48_Kernel43_Valid_Out, channel49_Kernel43_Valid_Out, channel50_Kernel43_Valid_Out, channel51_Kernel43_Valid_Out, channel52_Kernel43_Valid_Out, channel53_Kernel43_Valid_Out, channel54_Kernel43_Valid_Out, channel55_Kernel43_Valid_Out, channel56_Kernel43_Valid_Out, channel57_Kernel43_Valid_Out, channel58_Kernel43_Valid_Out, channel59_Kernel43_Valid_Out, channel60_Kernel43_Valid_Out, channel61_Kernel43_Valid_Out, channel62_Kernel43_Valid_Out, channel63_Kernel43_Valid_Out, channel64_Kernel43_Valid_Out;

	assign add_kernel43=channel1_Kernel43_Valid_Out & channel2_Kernel43_Valid_Out & channel3_Kernel43_Valid_Out & channel4_Kernel43_Valid_Out & channel5_Kernel43_Valid_Out & channel6_Kernel43_Valid_Out & channel7_Kernel43_Valid_Out & channel8_Kernel43_Valid_Out & channel9_Kernel43_Valid_Out & channel10_Kernel43_Valid_Out & channel11_Kernel43_Valid_Out & channel12_Kernel43_Valid_Out & channel13_Kernel43_Valid_Out & channel14_Kernel43_Valid_Out & channel15_Kernel43_Valid_Out & channel16_Kernel43_Valid_Out & channel17_Kernel43_Valid_Out & channel18_Kernel43_Valid_Out & channel19_Kernel43_Valid_Out & channel20_Kernel43_Valid_Out & channel21_Kernel43_Valid_Out & channel22_Kernel43_Valid_Out & channel23_Kernel43_Valid_Out & channel24_Kernel43_Valid_Out & channel25_Kernel43_Valid_Out & channel26_Kernel43_Valid_Out & channel27_Kernel43_Valid_Out & channel28_Kernel43_Valid_Out & channel29_Kernel43_Valid_Out & channel30_Kernel43_Valid_Out & channel31_Kernel43_Valid_Out & channel32_Kernel43_Valid_Out & channel33_Kernel43_Valid_Out & channel34_Kernel43_Valid_Out & channel35_Kernel43_Valid_Out & channel36_Kernel43_Valid_Out & channel37_Kernel43_Valid_Out & channel38_Kernel43_Valid_Out & channel39_Kernel43_Valid_Out & channel40_Kernel43_Valid_Out & channel41_Kernel43_Valid_Out & channel42_Kernel43_Valid_Out & channel43_Kernel43_Valid_Out & channel44_Kernel43_Valid_Out & channel45_Kernel43_Valid_Out & channel46_Kernel43_Valid_Out & channel47_Kernel43_Valid_Out & channel48_Kernel43_Valid_Out & channel49_Kernel43_Valid_Out & channel50_Kernel43_Valid_Out & channel51_Kernel43_Valid_Out & channel52_Kernel43_Valid_Out & channel53_Kernel43_Valid_Out & channel54_Kernel43_Valid_Out & channel55_Kernel43_Valid_Out & channel56_Kernel43_Valid_Out & channel57_Kernel43_Valid_Out & channel58_Kernel43_Valid_Out & channel59_Kernel43_Valid_Out & channel60_Kernel43_Valid_Out & channel61_Kernel43_Valid_Out & channel62_Kernel43_Valid_Out & channel63_Kernel43_Valid_Out & channel64_Kernel43_Valid_Out;

	wire channel1_Kernel44_Valid_Out, channel2_Kernel44_Valid_Out, channel3_Kernel44_Valid_Out, channel4_Kernel44_Valid_Out, channel5_Kernel44_Valid_Out, channel6_Kernel44_Valid_Out, channel7_Kernel44_Valid_Out, channel8_Kernel44_Valid_Out, channel9_Kernel44_Valid_Out, channel10_Kernel44_Valid_Out, channel11_Kernel44_Valid_Out, channel12_Kernel44_Valid_Out, channel13_Kernel44_Valid_Out, channel14_Kernel44_Valid_Out, channel15_Kernel44_Valid_Out, channel16_Kernel44_Valid_Out, channel17_Kernel44_Valid_Out, channel18_Kernel44_Valid_Out, channel19_Kernel44_Valid_Out, channel20_Kernel44_Valid_Out, channel21_Kernel44_Valid_Out, channel22_Kernel44_Valid_Out, channel23_Kernel44_Valid_Out, channel24_Kernel44_Valid_Out, channel25_Kernel44_Valid_Out, channel26_Kernel44_Valid_Out, channel27_Kernel44_Valid_Out, channel28_Kernel44_Valid_Out, channel29_Kernel44_Valid_Out, channel30_Kernel44_Valid_Out, channel31_Kernel44_Valid_Out, channel32_Kernel44_Valid_Out, channel33_Kernel44_Valid_Out, channel34_Kernel44_Valid_Out, channel35_Kernel44_Valid_Out, channel36_Kernel44_Valid_Out, channel37_Kernel44_Valid_Out, channel38_Kernel44_Valid_Out, channel39_Kernel44_Valid_Out, channel40_Kernel44_Valid_Out, channel41_Kernel44_Valid_Out, channel42_Kernel44_Valid_Out, channel43_Kernel44_Valid_Out, channel44_Kernel44_Valid_Out, channel45_Kernel44_Valid_Out, channel46_Kernel44_Valid_Out, channel47_Kernel44_Valid_Out, channel48_Kernel44_Valid_Out, channel49_Kernel44_Valid_Out, channel50_Kernel44_Valid_Out, channel51_Kernel44_Valid_Out, channel52_Kernel44_Valid_Out, channel53_Kernel44_Valid_Out, channel54_Kernel44_Valid_Out, channel55_Kernel44_Valid_Out, channel56_Kernel44_Valid_Out, channel57_Kernel44_Valid_Out, channel58_Kernel44_Valid_Out, channel59_Kernel44_Valid_Out, channel60_Kernel44_Valid_Out, channel61_Kernel44_Valid_Out, channel62_Kernel44_Valid_Out, channel63_Kernel44_Valid_Out, channel64_Kernel44_Valid_Out;

	assign add_kernel44=channel1_Kernel44_Valid_Out & channel2_Kernel44_Valid_Out & channel3_Kernel44_Valid_Out & channel4_Kernel44_Valid_Out & channel5_Kernel44_Valid_Out & channel6_Kernel44_Valid_Out & channel7_Kernel44_Valid_Out & channel8_Kernel44_Valid_Out & channel9_Kernel44_Valid_Out & channel10_Kernel44_Valid_Out & channel11_Kernel44_Valid_Out & channel12_Kernel44_Valid_Out & channel13_Kernel44_Valid_Out & channel14_Kernel44_Valid_Out & channel15_Kernel44_Valid_Out & channel16_Kernel44_Valid_Out & channel17_Kernel44_Valid_Out & channel18_Kernel44_Valid_Out & channel19_Kernel44_Valid_Out & channel20_Kernel44_Valid_Out & channel21_Kernel44_Valid_Out & channel22_Kernel44_Valid_Out & channel23_Kernel44_Valid_Out & channel24_Kernel44_Valid_Out & channel25_Kernel44_Valid_Out & channel26_Kernel44_Valid_Out & channel27_Kernel44_Valid_Out & channel28_Kernel44_Valid_Out & channel29_Kernel44_Valid_Out & channel30_Kernel44_Valid_Out & channel31_Kernel44_Valid_Out & channel32_Kernel44_Valid_Out & channel33_Kernel44_Valid_Out & channel34_Kernel44_Valid_Out & channel35_Kernel44_Valid_Out & channel36_Kernel44_Valid_Out & channel37_Kernel44_Valid_Out & channel38_Kernel44_Valid_Out & channel39_Kernel44_Valid_Out & channel40_Kernel44_Valid_Out & channel41_Kernel44_Valid_Out & channel42_Kernel44_Valid_Out & channel43_Kernel44_Valid_Out & channel44_Kernel44_Valid_Out & channel45_Kernel44_Valid_Out & channel46_Kernel44_Valid_Out & channel47_Kernel44_Valid_Out & channel48_Kernel44_Valid_Out & channel49_Kernel44_Valid_Out & channel50_Kernel44_Valid_Out & channel51_Kernel44_Valid_Out & channel52_Kernel44_Valid_Out & channel53_Kernel44_Valid_Out & channel54_Kernel44_Valid_Out & channel55_Kernel44_Valid_Out & channel56_Kernel44_Valid_Out & channel57_Kernel44_Valid_Out & channel58_Kernel44_Valid_Out & channel59_Kernel44_Valid_Out & channel60_Kernel44_Valid_Out & channel61_Kernel44_Valid_Out & channel62_Kernel44_Valid_Out & channel63_Kernel44_Valid_Out & channel64_Kernel44_Valid_Out;

	wire channel1_Kernel45_Valid_Out, channel2_Kernel45_Valid_Out, channel3_Kernel45_Valid_Out, channel4_Kernel45_Valid_Out, channel5_Kernel45_Valid_Out, channel6_Kernel45_Valid_Out, channel7_Kernel45_Valid_Out, channel8_Kernel45_Valid_Out, channel9_Kernel45_Valid_Out, channel10_Kernel45_Valid_Out, channel11_Kernel45_Valid_Out, channel12_Kernel45_Valid_Out, channel13_Kernel45_Valid_Out, channel14_Kernel45_Valid_Out, channel15_Kernel45_Valid_Out, channel16_Kernel45_Valid_Out, channel17_Kernel45_Valid_Out, channel18_Kernel45_Valid_Out, channel19_Kernel45_Valid_Out, channel20_Kernel45_Valid_Out, channel21_Kernel45_Valid_Out, channel22_Kernel45_Valid_Out, channel23_Kernel45_Valid_Out, channel24_Kernel45_Valid_Out, channel25_Kernel45_Valid_Out, channel26_Kernel45_Valid_Out, channel27_Kernel45_Valid_Out, channel28_Kernel45_Valid_Out, channel29_Kernel45_Valid_Out, channel30_Kernel45_Valid_Out, channel31_Kernel45_Valid_Out, channel32_Kernel45_Valid_Out, channel33_Kernel45_Valid_Out, channel34_Kernel45_Valid_Out, channel35_Kernel45_Valid_Out, channel36_Kernel45_Valid_Out, channel37_Kernel45_Valid_Out, channel38_Kernel45_Valid_Out, channel39_Kernel45_Valid_Out, channel40_Kernel45_Valid_Out, channel41_Kernel45_Valid_Out, channel42_Kernel45_Valid_Out, channel43_Kernel45_Valid_Out, channel44_Kernel45_Valid_Out, channel45_Kernel45_Valid_Out, channel46_Kernel45_Valid_Out, channel47_Kernel45_Valid_Out, channel48_Kernel45_Valid_Out, channel49_Kernel45_Valid_Out, channel50_Kernel45_Valid_Out, channel51_Kernel45_Valid_Out, channel52_Kernel45_Valid_Out, channel53_Kernel45_Valid_Out, channel54_Kernel45_Valid_Out, channel55_Kernel45_Valid_Out, channel56_Kernel45_Valid_Out, channel57_Kernel45_Valid_Out, channel58_Kernel45_Valid_Out, channel59_Kernel45_Valid_Out, channel60_Kernel45_Valid_Out, channel61_Kernel45_Valid_Out, channel62_Kernel45_Valid_Out, channel63_Kernel45_Valid_Out, channel64_Kernel45_Valid_Out;

	assign add_kernel45=channel1_Kernel45_Valid_Out & channel2_Kernel45_Valid_Out & channel3_Kernel45_Valid_Out & channel4_Kernel45_Valid_Out & channel5_Kernel45_Valid_Out & channel6_Kernel45_Valid_Out & channel7_Kernel45_Valid_Out & channel8_Kernel45_Valid_Out & channel9_Kernel45_Valid_Out & channel10_Kernel45_Valid_Out & channel11_Kernel45_Valid_Out & channel12_Kernel45_Valid_Out & channel13_Kernel45_Valid_Out & channel14_Kernel45_Valid_Out & channel15_Kernel45_Valid_Out & channel16_Kernel45_Valid_Out & channel17_Kernel45_Valid_Out & channel18_Kernel45_Valid_Out & channel19_Kernel45_Valid_Out & channel20_Kernel45_Valid_Out & channel21_Kernel45_Valid_Out & channel22_Kernel45_Valid_Out & channel23_Kernel45_Valid_Out & channel24_Kernel45_Valid_Out & channel25_Kernel45_Valid_Out & channel26_Kernel45_Valid_Out & channel27_Kernel45_Valid_Out & channel28_Kernel45_Valid_Out & channel29_Kernel45_Valid_Out & channel30_Kernel45_Valid_Out & channel31_Kernel45_Valid_Out & channel32_Kernel45_Valid_Out & channel33_Kernel45_Valid_Out & channel34_Kernel45_Valid_Out & channel35_Kernel45_Valid_Out & channel36_Kernel45_Valid_Out & channel37_Kernel45_Valid_Out & channel38_Kernel45_Valid_Out & channel39_Kernel45_Valid_Out & channel40_Kernel45_Valid_Out & channel41_Kernel45_Valid_Out & channel42_Kernel45_Valid_Out & channel43_Kernel45_Valid_Out & channel44_Kernel45_Valid_Out & channel45_Kernel45_Valid_Out & channel46_Kernel45_Valid_Out & channel47_Kernel45_Valid_Out & channel48_Kernel45_Valid_Out & channel49_Kernel45_Valid_Out & channel50_Kernel45_Valid_Out & channel51_Kernel45_Valid_Out & channel52_Kernel45_Valid_Out & channel53_Kernel45_Valid_Out & channel54_Kernel45_Valid_Out & channel55_Kernel45_Valid_Out & channel56_Kernel45_Valid_Out & channel57_Kernel45_Valid_Out & channel58_Kernel45_Valid_Out & channel59_Kernel45_Valid_Out & channel60_Kernel45_Valid_Out & channel61_Kernel45_Valid_Out & channel62_Kernel45_Valid_Out & channel63_Kernel45_Valid_Out & channel64_Kernel45_Valid_Out;

	wire channel1_Kernel46_Valid_Out, channel2_Kernel46_Valid_Out, channel3_Kernel46_Valid_Out, channel4_Kernel46_Valid_Out, channel5_Kernel46_Valid_Out, channel6_Kernel46_Valid_Out, channel7_Kernel46_Valid_Out, channel8_Kernel46_Valid_Out, channel9_Kernel46_Valid_Out, channel10_Kernel46_Valid_Out, channel11_Kernel46_Valid_Out, channel12_Kernel46_Valid_Out, channel13_Kernel46_Valid_Out, channel14_Kernel46_Valid_Out, channel15_Kernel46_Valid_Out, channel16_Kernel46_Valid_Out, channel17_Kernel46_Valid_Out, channel18_Kernel46_Valid_Out, channel19_Kernel46_Valid_Out, channel20_Kernel46_Valid_Out, channel21_Kernel46_Valid_Out, channel22_Kernel46_Valid_Out, channel23_Kernel46_Valid_Out, channel24_Kernel46_Valid_Out, channel25_Kernel46_Valid_Out, channel26_Kernel46_Valid_Out, channel27_Kernel46_Valid_Out, channel28_Kernel46_Valid_Out, channel29_Kernel46_Valid_Out, channel30_Kernel46_Valid_Out, channel31_Kernel46_Valid_Out, channel32_Kernel46_Valid_Out, channel33_Kernel46_Valid_Out, channel34_Kernel46_Valid_Out, channel35_Kernel46_Valid_Out, channel36_Kernel46_Valid_Out, channel37_Kernel46_Valid_Out, channel38_Kernel46_Valid_Out, channel39_Kernel46_Valid_Out, channel40_Kernel46_Valid_Out, channel41_Kernel46_Valid_Out, channel42_Kernel46_Valid_Out, channel43_Kernel46_Valid_Out, channel44_Kernel46_Valid_Out, channel45_Kernel46_Valid_Out, channel46_Kernel46_Valid_Out, channel47_Kernel46_Valid_Out, channel48_Kernel46_Valid_Out, channel49_Kernel46_Valid_Out, channel50_Kernel46_Valid_Out, channel51_Kernel46_Valid_Out, channel52_Kernel46_Valid_Out, channel53_Kernel46_Valid_Out, channel54_Kernel46_Valid_Out, channel55_Kernel46_Valid_Out, channel56_Kernel46_Valid_Out, channel57_Kernel46_Valid_Out, channel58_Kernel46_Valid_Out, channel59_Kernel46_Valid_Out, channel60_Kernel46_Valid_Out, channel61_Kernel46_Valid_Out, channel62_Kernel46_Valid_Out, channel63_Kernel46_Valid_Out, channel64_Kernel46_Valid_Out;

	assign add_kernel46=channel1_Kernel46_Valid_Out & channel2_Kernel46_Valid_Out & channel3_Kernel46_Valid_Out & channel4_Kernel46_Valid_Out & channel5_Kernel46_Valid_Out & channel6_Kernel46_Valid_Out & channel7_Kernel46_Valid_Out & channel8_Kernel46_Valid_Out & channel9_Kernel46_Valid_Out & channel10_Kernel46_Valid_Out & channel11_Kernel46_Valid_Out & channel12_Kernel46_Valid_Out & channel13_Kernel46_Valid_Out & channel14_Kernel46_Valid_Out & channel15_Kernel46_Valid_Out & channel16_Kernel46_Valid_Out & channel17_Kernel46_Valid_Out & channel18_Kernel46_Valid_Out & channel19_Kernel46_Valid_Out & channel20_Kernel46_Valid_Out & channel21_Kernel46_Valid_Out & channel22_Kernel46_Valid_Out & channel23_Kernel46_Valid_Out & channel24_Kernel46_Valid_Out & channel25_Kernel46_Valid_Out & channel26_Kernel46_Valid_Out & channel27_Kernel46_Valid_Out & channel28_Kernel46_Valid_Out & channel29_Kernel46_Valid_Out & channel30_Kernel46_Valid_Out & channel31_Kernel46_Valid_Out & channel32_Kernel46_Valid_Out & channel33_Kernel46_Valid_Out & channel34_Kernel46_Valid_Out & channel35_Kernel46_Valid_Out & channel36_Kernel46_Valid_Out & channel37_Kernel46_Valid_Out & channel38_Kernel46_Valid_Out & channel39_Kernel46_Valid_Out & channel40_Kernel46_Valid_Out & channel41_Kernel46_Valid_Out & channel42_Kernel46_Valid_Out & channel43_Kernel46_Valid_Out & channel44_Kernel46_Valid_Out & channel45_Kernel46_Valid_Out & channel46_Kernel46_Valid_Out & channel47_Kernel46_Valid_Out & channel48_Kernel46_Valid_Out & channel49_Kernel46_Valid_Out & channel50_Kernel46_Valid_Out & channel51_Kernel46_Valid_Out & channel52_Kernel46_Valid_Out & channel53_Kernel46_Valid_Out & channel54_Kernel46_Valid_Out & channel55_Kernel46_Valid_Out & channel56_Kernel46_Valid_Out & channel57_Kernel46_Valid_Out & channel58_Kernel46_Valid_Out & channel59_Kernel46_Valid_Out & channel60_Kernel46_Valid_Out & channel61_Kernel46_Valid_Out & channel62_Kernel46_Valid_Out & channel63_Kernel46_Valid_Out & channel64_Kernel46_Valid_Out;

	wire channel1_Kernel47_Valid_Out, channel2_Kernel47_Valid_Out, channel3_Kernel47_Valid_Out, channel4_Kernel47_Valid_Out, channel5_Kernel47_Valid_Out, channel6_Kernel47_Valid_Out, channel7_Kernel47_Valid_Out, channel8_Kernel47_Valid_Out, channel9_Kernel47_Valid_Out, channel10_Kernel47_Valid_Out, channel11_Kernel47_Valid_Out, channel12_Kernel47_Valid_Out, channel13_Kernel47_Valid_Out, channel14_Kernel47_Valid_Out, channel15_Kernel47_Valid_Out, channel16_Kernel47_Valid_Out, channel17_Kernel47_Valid_Out, channel18_Kernel47_Valid_Out, channel19_Kernel47_Valid_Out, channel20_Kernel47_Valid_Out, channel21_Kernel47_Valid_Out, channel22_Kernel47_Valid_Out, channel23_Kernel47_Valid_Out, channel24_Kernel47_Valid_Out, channel25_Kernel47_Valid_Out, channel26_Kernel47_Valid_Out, channel27_Kernel47_Valid_Out, channel28_Kernel47_Valid_Out, channel29_Kernel47_Valid_Out, channel30_Kernel47_Valid_Out, channel31_Kernel47_Valid_Out, channel32_Kernel47_Valid_Out, channel33_Kernel47_Valid_Out, channel34_Kernel47_Valid_Out, channel35_Kernel47_Valid_Out, channel36_Kernel47_Valid_Out, channel37_Kernel47_Valid_Out, channel38_Kernel47_Valid_Out, channel39_Kernel47_Valid_Out, channel40_Kernel47_Valid_Out, channel41_Kernel47_Valid_Out, channel42_Kernel47_Valid_Out, channel43_Kernel47_Valid_Out, channel44_Kernel47_Valid_Out, channel45_Kernel47_Valid_Out, channel46_Kernel47_Valid_Out, channel47_Kernel47_Valid_Out, channel48_Kernel47_Valid_Out, channel49_Kernel47_Valid_Out, channel50_Kernel47_Valid_Out, channel51_Kernel47_Valid_Out, channel52_Kernel47_Valid_Out, channel53_Kernel47_Valid_Out, channel54_Kernel47_Valid_Out, channel55_Kernel47_Valid_Out, channel56_Kernel47_Valid_Out, channel57_Kernel47_Valid_Out, channel58_Kernel47_Valid_Out, channel59_Kernel47_Valid_Out, channel60_Kernel47_Valid_Out, channel61_Kernel47_Valid_Out, channel62_Kernel47_Valid_Out, channel63_Kernel47_Valid_Out, channel64_Kernel47_Valid_Out;

	assign add_kernel47=channel1_Kernel47_Valid_Out & channel2_Kernel47_Valid_Out & channel3_Kernel47_Valid_Out & channel4_Kernel47_Valid_Out & channel5_Kernel47_Valid_Out & channel6_Kernel47_Valid_Out & channel7_Kernel47_Valid_Out & channel8_Kernel47_Valid_Out & channel9_Kernel47_Valid_Out & channel10_Kernel47_Valid_Out & channel11_Kernel47_Valid_Out & channel12_Kernel47_Valid_Out & channel13_Kernel47_Valid_Out & channel14_Kernel47_Valid_Out & channel15_Kernel47_Valid_Out & channel16_Kernel47_Valid_Out & channel17_Kernel47_Valid_Out & channel18_Kernel47_Valid_Out & channel19_Kernel47_Valid_Out & channel20_Kernel47_Valid_Out & channel21_Kernel47_Valid_Out & channel22_Kernel47_Valid_Out & channel23_Kernel47_Valid_Out & channel24_Kernel47_Valid_Out & channel25_Kernel47_Valid_Out & channel26_Kernel47_Valid_Out & channel27_Kernel47_Valid_Out & channel28_Kernel47_Valid_Out & channel29_Kernel47_Valid_Out & channel30_Kernel47_Valid_Out & channel31_Kernel47_Valid_Out & channel32_Kernel47_Valid_Out & channel33_Kernel47_Valid_Out & channel34_Kernel47_Valid_Out & channel35_Kernel47_Valid_Out & channel36_Kernel47_Valid_Out & channel37_Kernel47_Valid_Out & channel38_Kernel47_Valid_Out & channel39_Kernel47_Valid_Out & channel40_Kernel47_Valid_Out & channel41_Kernel47_Valid_Out & channel42_Kernel47_Valid_Out & channel43_Kernel47_Valid_Out & channel44_Kernel47_Valid_Out & channel45_Kernel47_Valid_Out & channel46_Kernel47_Valid_Out & channel47_Kernel47_Valid_Out & channel48_Kernel47_Valid_Out & channel49_Kernel47_Valid_Out & channel50_Kernel47_Valid_Out & channel51_Kernel47_Valid_Out & channel52_Kernel47_Valid_Out & channel53_Kernel47_Valid_Out & channel54_Kernel47_Valid_Out & channel55_Kernel47_Valid_Out & channel56_Kernel47_Valid_Out & channel57_Kernel47_Valid_Out & channel58_Kernel47_Valid_Out & channel59_Kernel47_Valid_Out & channel60_Kernel47_Valid_Out & channel61_Kernel47_Valid_Out & channel62_Kernel47_Valid_Out & channel63_Kernel47_Valid_Out & channel64_Kernel47_Valid_Out;

	wire channel1_Kernel48_Valid_Out, channel2_Kernel48_Valid_Out, channel3_Kernel48_Valid_Out, channel4_Kernel48_Valid_Out, channel5_Kernel48_Valid_Out, channel6_Kernel48_Valid_Out, channel7_Kernel48_Valid_Out, channel8_Kernel48_Valid_Out, channel9_Kernel48_Valid_Out, channel10_Kernel48_Valid_Out, channel11_Kernel48_Valid_Out, channel12_Kernel48_Valid_Out, channel13_Kernel48_Valid_Out, channel14_Kernel48_Valid_Out, channel15_Kernel48_Valid_Out, channel16_Kernel48_Valid_Out, channel17_Kernel48_Valid_Out, channel18_Kernel48_Valid_Out, channel19_Kernel48_Valid_Out, channel20_Kernel48_Valid_Out, channel21_Kernel48_Valid_Out, channel22_Kernel48_Valid_Out, channel23_Kernel48_Valid_Out, channel24_Kernel48_Valid_Out, channel25_Kernel48_Valid_Out, channel26_Kernel48_Valid_Out, channel27_Kernel48_Valid_Out, channel28_Kernel48_Valid_Out, channel29_Kernel48_Valid_Out, channel30_Kernel48_Valid_Out, channel31_Kernel48_Valid_Out, channel32_Kernel48_Valid_Out, channel33_Kernel48_Valid_Out, channel34_Kernel48_Valid_Out, channel35_Kernel48_Valid_Out, channel36_Kernel48_Valid_Out, channel37_Kernel48_Valid_Out, channel38_Kernel48_Valid_Out, channel39_Kernel48_Valid_Out, channel40_Kernel48_Valid_Out, channel41_Kernel48_Valid_Out, channel42_Kernel48_Valid_Out, channel43_Kernel48_Valid_Out, channel44_Kernel48_Valid_Out, channel45_Kernel48_Valid_Out, channel46_Kernel48_Valid_Out, channel47_Kernel48_Valid_Out, channel48_Kernel48_Valid_Out, channel49_Kernel48_Valid_Out, channel50_Kernel48_Valid_Out, channel51_Kernel48_Valid_Out, channel52_Kernel48_Valid_Out, channel53_Kernel48_Valid_Out, channel54_Kernel48_Valid_Out, channel55_Kernel48_Valid_Out, channel56_Kernel48_Valid_Out, channel57_Kernel48_Valid_Out, channel58_Kernel48_Valid_Out, channel59_Kernel48_Valid_Out, channel60_Kernel48_Valid_Out, channel61_Kernel48_Valid_Out, channel62_Kernel48_Valid_Out, channel63_Kernel48_Valid_Out, channel64_Kernel48_Valid_Out;

	assign add_kernel48=channel1_Kernel48_Valid_Out & channel2_Kernel48_Valid_Out & channel3_Kernel48_Valid_Out & channel4_Kernel48_Valid_Out & channel5_Kernel48_Valid_Out & channel6_Kernel48_Valid_Out & channel7_Kernel48_Valid_Out & channel8_Kernel48_Valid_Out & channel9_Kernel48_Valid_Out & channel10_Kernel48_Valid_Out & channel11_Kernel48_Valid_Out & channel12_Kernel48_Valid_Out & channel13_Kernel48_Valid_Out & channel14_Kernel48_Valid_Out & channel15_Kernel48_Valid_Out & channel16_Kernel48_Valid_Out & channel17_Kernel48_Valid_Out & channel18_Kernel48_Valid_Out & channel19_Kernel48_Valid_Out & channel20_Kernel48_Valid_Out & channel21_Kernel48_Valid_Out & channel22_Kernel48_Valid_Out & channel23_Kernel48_Valid_Out & channel24_Kernel48_Valid_Out & channel25_Kernel48_Valid_Out & channel26_Kernel48_Valid_Out & channel27_Kernel48_Valid_Out & channel28_Kernel48_Valid_Out & channel29_Kernel48_Valid_Out & channel30_Kernel48_Valid_Out & channel31_Kernel48_Valid_Out & channel32_Kernel48_Valid_Out & channel33_Kernel48_Valid_Out & channel34_Kernel48_Valid_Out & channel35_Kernel48_Valid_Out & channel36_Kernel48_Valid_Out & channel37_Kernel48_Valid_Out & channel38_Kernel48_Valid_Out & channel39_Kernel48_Valid_Out & channel40_Kernel48_Valid_Out & channel41_Kernel48_Valid_Out & channel42_Kernel48_Valid_Out & channel43_Kernel48_Valid_Out & channel44_Kernel48_Valid_Out & channel45_Kernel48_Valid_Out & channel46_Kernel48_Valid_Out & channel47_Kernel48_Valid_Out & channel48_Kernel48_Valid_Out & channel49_Kernel48_Valid_Out & channel50_Kernel48_Valid_Out & channel51_Kernel48_Valid_Out & channel52_Kernel48_Valid_Out & channel53_Kernel48_Valid_Out & channel54_Kernel48_Valid_Out & channel55_Kernel48_Valid_Out & channel56_Kernel48_Valid_Out & channel57_Kernel48_Valid_Out & channel58_Kernel48_Valid_Out & channel59_Kernel48_Valid_Out & channel60_Kernel48_Valid_Out & channel61_Kernel48_Valid_Out & channel62_Kernel48_Valid_Out & channel63_Kernel48_Valid_Out & channel64_Kernel48_Valid_Out;

	wire channel1_Kernel49_Valid_Out, channel2_Kernel49_Valid_Out, channel3_Kernel49_Valid_Out, channel4_Kernel49_Valid_Out, channel5_Kernel49_Valid_Out, channel6_Kernel49_Valid_Out, channel7_Kernel49_Valid_Out, channel8_Kernel49_Valid_Out, channel9_Kernel49_Valid_Out, channel10_Kernel49_Valid_Out, channel11_Kernel49_Valid_Out, channel12_Kernel49_Valid_Out, channel13_Kernel49_Valid_Out, channel14_Kernel49_Valid_Out, channel15_Kernel49_Valid_Out, channel16_Kernel49_Valid_Out, channel17_Kernel49_Valid_Out, channel18_Kernel49_Valid_Out, channel19_Kernel49_Valid_Out, channel20_Kernel49_Valid_Out, channel21_Kernel49_Valid_Out, channel22_Kernel49_Valid_Out, channel23_Kernel49_Valid_Out, channel24_Kernel49_Valid_Out, channel25_Kernel49_Valid_Out, channel26_Kernel49_Valid_Out, channel27_Kernel49_Valid_Out, channel28_Kernel49_Valid_Out, channel29_Kernel49_Valid_Out, channel30_Kernel49_Valid_Out, channel31_Kernel49_Valid_Out, channel32_Kernel49_Valid_Out, channel33_Kernel49_Valid_Out, channel34_Kernel49_Valid_Out, channel35_Kernel49_Valid_Out, channel36_Kernel49_Valid_Out, channel37_Kernel49_Valid_Out, channel38_Kernel49_Valid_Out, channel39_Kernel49_Valid_Out, channel40_Kernel49_Valid_Out, channel41_Kernel49_Valid_Out, channel42_Kernel49_Valid_Out, channel43_Kernel49_Valid_Out, channel44_Kernel49_Valid_Out, channel45_Kernel49_Valid_Out, channel46_Kernel49_Valid_Out, channel47_Kernel49_Valid_Out, channel48_Kernel49_Valid_Out, channel49_Kernel49_Valid_Out, channel50_Kernel49_Valid_Out, channel51_Kernel49_Valid_Out, channel52_Kernel49_Valid_Out, channel53_Kernel49_Valid_Out, channel54_Kernel49_Valid_Out, channel55_Kernel49_Valid_Out, channel56_Kernel49_Valid_Out, channel57_Kernel49_Valid_Out, channel58_Kernel49_Valid_Out, channel59_Kernel49_Valid_Out, channel60_Kernel49_Valid_Out, channel61_Kernel49_Valid_Out, channel62_Kernel49_Valid_Out, channel63_Kernel49_Valid_Out, channel64_Kernel49_Valid_Out;

	assign add_kernel49=channel1_Kernel49_Valid_Out & channel2_Kernel49_Valid_Out & channel3_Kernel49_Valid_Out & channel4_Kernel49_Valid_Out & channel5_Kernel49_Valid_Out & channel6_Kernel49_Valid_Out & channel7_Kernel49_Valid_Out & channel8_Kernel49_Valid_Out & channel9_Kernel49_Valid_Out & channel10_Kernel49_Valid_Out & channel11_Kernel49_Valid_Out & channel12_Kernel49_Valid_Out & channel13_Kernel49_Valid_Out & channel14_Kernel49_Valid_Out & channel15_Kernel49_Valid_Out & channel16_Kernel49_Valid_Out & channel17_Kernel49_Valid_Out & channel18_Kernel49_Valid_Out & channel19_Kernel49_Valid_Out & channel20_Kernel49_Valid_Out & channel21_Kernel49_Valid_Out & channel22_Kernel49_Valid_Out & channel23_Kernel49_Valid_Out & channel24_Kernel49_Valid_Out & channel25_Kernel49_Valid_Out & channel26_Kernel49_Valid_Out & channel27_Kernel49_Valid_Out & channel28_Kernel49_Valid_Out & channel29_Kernel49_Valid_Out & channel30_Kernel49_Valid_Out & channel31_Kernel49_Valid_Out & channel32_Kernel49_Valid_Out & channel33_Kernel49_Valid_Out & channel34_Kernel49_Valid_Out & channel35_Kernel49_Valid_Out & channel36_Kernel49_Valid_Out & channel37_Kernel49_Valid_Out & channel38_Kernel49_Valid_Out & channel39_Kernel49_Valid_Out & channel40_Kernel49_Valid_Out & channel41_Kernel49_Valid_Out & channel42_Kernel49_Valid_Out & channel43_Kernel49_Valid_Out & channel44_Kernel49_Valid_Out & channel45_Kernel49_Valid_Out & channel46_Kernel49_Valid_Out & channel47_Kernel49_Valid_Out & channel48_Kernel49_Valid_Out & channel49_Kernel49_Valid_Out & channel50_Kernel49_Valid_Out & channel51_Kernel49_Valid_Out & channel52_Kernel49_Valid_Out & channel53_Kernel49_Valid_Out & channel54_Kernel49_Valid_Out & channel55_Kernel49_Valid_Out & channel56_Kernel49_Valid_Out & channel57_Kernel49_Valid_Out & channel58_Kernel49_Valid_Out & channel59_Kernel49_Valid_Out & channel60_Kernel49_Valid_Out & channel61_Kernel49_Valid_Out & channel62_Kernel49_Valid_Out & channel63_Kernel49_Valid_Out & channel64_Kernel49_Valid_Out;

	wire channel1_Kernel50_Valid_Out, channel2_Kernel50_Valid_Out, channel3_Kernel50_Valid_Out, channel4_Kernel50_Valid_Out, channel5_Kernel50_Valid_Out, channel6_Kernel50_Valid_Out, channel7_Kernel50_Valid_Out, channel8_Kernel50_Valid_Out, channel9_Kernel50_Valid_Out, channel10_Kernel50_Valid_Out, channel11_Kernel50_Valid_Out, channel12_Kernel50_Valid_Out, channel13_Kernel50_Valid_Out, channel14_Kernel50_Valid_Out, channel15_Kernel50_Valid_Out, channel16_Kernel50_Valid_Out, channel17_Kernel50_Valid_Out, channel18_Kernel50_Valid_Out, channel19_Kernel50_Valid_Out, channel20_Kernel50_Valid_Out, channel21_Kernel50_Valid_Out, channel22_Kernel50_Valid_Out, channel23_Kernel50_Valid_Out, channel24_Kernel50_Valid_Out, channel25_Kernel50_Valid_Out, channel26_Kernel50_Valid_Out, channel27_Kernel50_Valid_Out, channel28_Kernel50_Valid_Out, channel29_Kernel50_Valid_Out, channel30_Kernel50_Valid_Out, channel31_Kernel50_Valid_Out, channel32_Kernel50_Valid_Out, channel33_Kernel50_Valid_Out, channel34_Kernel50_Valid_Out, channel35_Kernel50_Valid_Out, channel36_Kernel50_Valid_Out, channel37_Kernel50_Valid_Out, channel38_Kernel50_Valid_Out, channel39_Kernel50_Valid_Out, channel40_Kernel50_Valid_Out, channel41_Kernel50_Valid_Out, channel42_Kernel50_Valid_Out, channel43_Kernel50_Valid_Out, channel44_Kernel50_Valid_Out, channel45_Kernel50_Valid_Out, channel46_Kernel50_Valid_Out, channel47_Kernel50_Valid_Out, channel48_Kernel50_Valid_Out, channel49_Kernel50_Valid_Out, channel50_Kernel50_Valid_Out, channel51_Kernel50_Valid_Out, channel52_Kernel50_Valid_Out, channel53_Kernel50_Valid_Out, channel54_Kernel50_Valid_Out, channel55_Kernel50_Valid_Out, channel56_Kernel50_Valid_Out, channel57_Kernel50_Valid_Out, channel58_Kernel50_Valid_Out, channel59_Kernel50_Valid_Out, channel60_Kernel50_Valid_Out, channel61_Kernel50_Valid_Out, channel62_Kernel50_Valid_Out, channel63_Kernel50_Valid_Out, channel64_Kernel50_Valid_Out;

	assign add_kernel50=channel1_Kernel50_Valid_Out & channel2_Kernel50_Valid_Out & channel3_Kernel50_Valid_Out & channel4_Kernel50_Valid_Out & channel5_Kernel50_Valid_Out & channel6_Kernel50_Valid_Out & channel7_Kernel50_Valid_Out & channel8_Kernel50_Valid_Out & channel9_Kernel50_Valid_Out & channel10_Kernel50_Valid_Out & channel11_Kernel50_Valid_Out & channel12_Kernel50_Valid_Out & channel13_Kernel50_Valid_Out & channel14_Kernel50_Valid_Out & channel15_Kernel50_Valid_Out & channel16_Kernel50_Valid_Out & channel17_Kernel50_Valid_Out & channel18_Kernel50_Valid_Out & channel19_Kernel50_Valid_Out & channel20_Kernel50_Valid_Out & channel21_Kernel50_Valid_Out & channel22_Kernel50_Valid_Out & channel23_Kernel50_Valid_Out & channel24_Kernel50_Valid_Out & channel25_Kernel50_Valid_Out & channel26_Kernel50_Valid_Out & channel27_Kernel50_Valid_Out & channel28_Kernel50_Valid_Out & channel29_Kernel50_Valid_Out & channel30_Kernel50_Valid_Out & channel31_Kernel50_Valid_Out & channel32_Kernel50_Valid_Out & channel33_Kernel50_Valid_Out & channel34_Kernel50_Valid_Out & channel35_Kernel50_Valid_Out & channel36_Kernel50_Valid_Out & channel37_Kernel50_Valid_Out & channel38_Kernel50_Valid_Out & channel39_Kernel50_Valid_Out & channel40_Kernel50_Valid_Out & channel41_Kernel50_Valid_Out & channel42_Kernel50_Valid_Out & channel43_Kernel50_Valid_Out & channel44_Kernel50_Valid_Out & channel45_Kernel50_Valid_Out & channel46_Kernel50_Valid_Out & channel47_Kernel50_Valid_Out & channel48_Kernel50_Valid_Out & channel49_Kernel50_Valid_Out & channel50_Kernel50_Valid_Out & channel51_Kernel50_Valid_Out & channel52_Kernel50_Valid_Out & channel53_Kernel50_Valid_Out & channel54_Kernel50_Valid_Out & channel55_Kernel50_Valid_Out & channel56_Kernel50_Valid_Out & channel57_Kernel50_Valid_Out & channel58_Kernel50_Valid_Out & channel59_Kernel50_Valid_Out & channel60_Kernel50_Valid_Out & channel61_Kernel50_Valid_Out & channel62_Kernel50_Valid_Out & channel63_Kernel50_Valid_Out & channel64_Kernel50_Valid_Out;

	wire channel1_Kernel51_Valid_Out, channel2_Kernel51_Valid_Out, channel3_Kernel51_Valid_Out, channel4_Kernel51_Valid_Out, channel5_Kernel51_Valid_Out, channel6_Kernel51_Valid_Out, channel7_Kernel51_Valid_Out, channel8_Kernel51_Valid_Out, channel9_Kernel51_Valid_Out, channel10_Kernel51_Valid_Out, channel11_Kernel51_Valid_Out, channel12_Kernel51_Valid_Out, channel13_Kernel51_Valid_Out, channel14_Kernel51_Valid_Out, channel15_Kernel51_Valid_Out, channel16_Kernel51_Valid_Out, channel17_Kernel51_Valid_Out, channel18_Kernel51_Valid_Out, channel19_Kernel51_Valid_Out, channel20_Kernel51_Valid_Out, channel21_Kernel51_Valid_Out, channel22_Kernel51_Valid_Out, channel23_Kernel51_Valid_Out, channel24_Kernel51_Valid_Out, channel25_Kernel51_Valid_Out, channel26_Kernel51_Valid_Out, channel27_Kernel51_Valid_Out, channel28_Kernel51_Valid_Out, channel29_Kernel51_Valid_Out, channel30_Kernel51_Valid_Out, channel31_Kernel51_Valid_Out, channel32_Kernel51_Valid_Out, channel33_Kernel51_Valid_Out, channel34_Kernel51_Valid_Out, channel35_Kernel51_Valid_Out, channel36_Kernel51_Valid_Out, channel37_Kernel51_Valid_Out, channel38_Kernel51_Valid_Out, channel39_Kernel51_Valid_Out, channel40_Kernel51_Valid_Out, channel41_Kernel51_Valid_Out, channel42_Kernel51_Valid_Out, channel43_Kernel51_Valid_Out, channel44_Kernel51_Valid_Out, channel45_Kernel51_Valid_Out, channel46_Kernel51_Valid_Out, channel47_Kernel51_Valid_Out, channel48_Kernel51_Valid_Out, channel49_Kernel51_Valid_Out, channel50_Kernel51_Valid_Out, channel51_Kernel51_Valid_Out, channel52_Kernel51_Valid_Out, channel53_Kernel51_Valid_Out, channel54_Kernel51_Valid_Out, channel55_Kernel51_Valid_Out, channel56_Kernel51_Valid_Out, channel57_Kernel51_Valid_Out, channel58_Kernel51_Valid_Out, channel59_Kernel51_Valid_Out, channel60_Kernel51_Valid_Out, channel61_Kernel51_Valid_Out, channel62_Kernel51_Valid_Out, channel63_Kernel51_Valid_Out, channel64_Kernel51_Valid_Out;

	assign add_kernel51=channel1_Kernel51_Valid_Out & channel2_Kernel51_Valid_Out & channel3_Kernel51_Valid_Out & channel4_Kernel51_Valid_Out & channel5_Kernel51_Valid_Out & channel6_Kernel51_Valid_Out & channel7_Kernel51_Valid_Out & channel8_Kernel51_Valid_Out & channel9_Kernel51_Valid_Out & channel10_Kernel51_Valid_Out & channel11_Kernel51_Valid_Out & channel12_Kernel51_Valid_Out & channel13_Kernel51_Valid_Out & channel14_Kernel51_Valid_Out & channel15_Kernel51_Valid_Out & channel16_Kernel51_Valid_Out & channel17_Kernel51_Valid_Out & channel18_Kernel51_Valid_Out & channel19_Kernel51_Valid_Out & channel20_Kernel51_Valid_Out & channel21_Kernel51_Valid_Out & channel22_Kernel51_Valid_Out & channel23_Kernel51_Valid_Out & channel24_Kernel51_Valid_Out & channel25_Kernel51_Valid_Out & channel26_Kernel51_Valid_Out & channel27_Kernel51_Valid_Out & channel28_Kernel51_Valid_Out & channel29_Kernel51_Valid_Out & channel30_Kernel51_Valid_Out & channel31_Kernel51_Valid_Out & channel32_Kernel51_Valid_Out & channel33_Kernel51_Valid_Out & channel34_Kernel51_Valid_Out & channel35_Kernel51_Valid_Out & channel36_Kernel51_Valid_Out & channel37_Kernel51_Valid_Out & channel38_Kernel51_Valid_Out & channel39_Kernel51_Valid_Out & channel40_Kernel51_Valid_Out & channel41_Kernel51_Valid_Out & channel42_Kernel51_Valid_Out & channel43_Kernel51_Valid_Out & channel44_Kernel51_Valid_Out & channel45_Kernel51_Valid_Out & channel46_Kernel51_Valid_Out & channel47_Kernel51_Valid_Out & channel48_Kernel51_Valid_Out & channel49_Kernel51_Valid_Out & channel50_Kernel51_Valid_Out & channel51_Kernel51_Valid_Out & channel52_Kernel51_Valid_Out & channel53_Kernel51_Valid_Out & channel54_Kernel51_Valid_Out & channel55_Kernel51_Valid_Out & channel56_Kernel51_Valid_Out & channel57_Kernel51_Valid_Out & channel58_Kernel51_Valid_Out & channel59_Kernel51_Valid_Out & channel60_Kernel51_Valid_Out & channel61_Kernel51_Valid_Out & channel62_Kernel51_Valid_Out & channel63_Kernel51_Valid_Out & channel64_Kernel51_Valid_Out;

	wire channel1_Kernel52_Valid_Out, channel2_Kernel52_Valid_Out, channel3_Kernel52_Valid_Out, channel4_Kernel52_Valid_Out, channel5_Kernel52_Valid_Out, channel6_Kernel52_Valid_Out, channel7_Kernel52_Valid_Out, channel8_Kernel52_Valid_Out, channel9_Kernel52_Valid_Out, channel10_Kernel52_Valid_Out, channel11_Kernel52_Valid_Out, channel12_Kernel52_Valid_Out, channel13_Kernel52_Valid_Out, channel14_Kernel52_Valid_Out, channel15_Kernel52_Valid_Out, channel16_Kernel52_Valid_Out, channel17_Kernel52_Valid_Out, channel18_Kernel52_Valid_Out, channel19_Kernel52_Valid_Out, channel20_Kernel52_Valid_Out, channel21_Kernel52_Valid_Out, channel22_Kernel52_Valid_Out, channel23_Kernel52_Valid_Out, channel24_Kernel52_Valid_Out, channel25_Kernel52_Valid_Out, channel26_Kernel52_Valid_Out, channel27_Kernel52_Valid_Out, channel28_Kernel52_Valid_Out, channel29_Kernel52_Valid_Out, channel30_Kernel52_Valid_Out, channel31_Kernel52_Valid_Out, channel32_Kernel52_Valid_Out, channel33_Kernel52_Valid_Out, channel34_Kernel52_Valid_Out, channel35_Kernel52_Valid_Out, channel36_Kernel52_Valid_Out, channel37_Kernel52_Valid_Out, channel38_Kernel52_Valid_Out, channel39_Kernel52_Valid_Out, channel40_Kernel52_Valid_Out, channel41_Kernel52_Valid_Out, channel42_Kernel52_Valid_Out, channel43_Kernel52_Valid_Out, channel44_Kernel52_Valid_Out, channel45_Kernel52_Valid_Out, channel46_Kernel52_Valid_Out, channel47_Kernel52_Valid_Out, channel48_Kernel52_Valid_Out, channel49_Kernel52_Valid_Out, channel50_Kernel52_Valid_Out, channel51_Kernel52_Valid_Out, channel52_Kernel52_Valid_Out, channel53_Kernel52_Valid_Out, channel54_Kernel52_Valid_Out, channel55_Kernel52_Valid_Out, channel56_Kernel52_Valid_Out, channel57_Kernel52_Valid_Out, channel58_Kernel52_Valid_Out, channel59_Kernel52_Valid_Out, channel60_Kernel52_Valid_Out, channel61_Kernel52_Valid_Out, channel62_Kernel52_Valid_Out, channel63_Kernel52_Valid_Out, channel64_Kernel52_Valid_Out;

	assign add_kernel52=channel1_Kernel52_Valid_Out & channel2_Kernel52_Valid_Out & channel3_Kernel52_Valid_Out & channel4_Kernel52_Valid_Out & channel5_Kernel52_Valid_Out & channel6_Kernel52_Valid_Out & channel7_Kernel52_Valid_Out & channel8_Kernel52_Valid_Out & channel9_Kernel52_Valid_Out & channel10_Kernel52_Valid_Out & channel11_Kernel52_Valid_Out & channel12_Kernel52_Valid_Out & channel13_Kernel52_Valid_Out & channel14_Kernel52_Valid_Out & channel15_Kernel52_Valid_Out & channel16_Kernel52_Valid_Out & channel17_Kernel52_Valid_Out & channel18_Kernel52_Valid_Out & channel19_Kernel52_Valid_Out & channel20_Kernel52_Valid_Out & channel21_Kernel52_Valid_Out & channel22_Kernel52_Valid_Out & channel23_Kernel52_Valid_Out & channel24_Kernel52_Valid_Out & channel25_Kernel52_Valid_Out & channel26_Kernel52_Valid_Out & channel27_Kernel52_Valid_Out & channel28_Kernel52_Valid_Out & channel29_Kernel52_Valid_Out & channel30_Kernel52_Valid_Out & channel31_Kernel52_Valid_Out & channel32_Kernel52_Valid_Out & channel33_Kernel52_Valid_Out & channel34_Kernel52_Valid_Out & channel35_Kernel52_Valid_Out & channel36_Kernel52_Valid_Out & channel37_Kernel52_Valid_Out & channel38_Kernel52_Valid_Out & channel39_Kernel52_Valid_Out & channel40_Kernel52_Valid_Out & channel41_Kernel52_Valid_Out & channel42_Kernel52_Valid_Out & channel43_Kernel52_Valid_Out & channel44_Kernel52_Valid_Out & channel45_Kernel52_Valid_Out & channel46_Kernel52_Valid_Out & channel47_Kernel52_Valid_Out & channel48_Kernel52_Valid_Out & channel49_Kernel52_Valid_Out & channel50_Kernel52_Valid_Out & channel51_Kernel52_Valid_Out & channel52_Kernel52_Valid_Out & channel53_Kernel52_Valid_Out & channel54_Kernel52_Valid_Out & channel55_Kernel52_Valid_Out & channel56_Kernel52_Valid_Out & channel57_Kernel52_Valid_Out & channel58_Kernel52_Valid_Out & channel59_Kernel52_Valid_Out & channel60_Kernel52_Valid_Out & channel61_Kernel52_Valid_Out & channel62_Kernel52_Valid_Out & channel63_Kernel52_Valid_Out & channel64_Kernel52_Valid_Out;

	wire channel1_Kernel53_Valid_Out, channel2_Kernel53_Valid_Out, channel3_Kernel53_Valid_Out, channel4_Kernel53_Valid_Out, channel5_Kernel53_Valid_Out, channel6_Kernel53_Valid_Out, channel7_Kernel53_Valid_Out, channel8_Kernel53_Valid_Out, channel9_Kernel53_Valid_Out, channel10_Kernel53_Valid_Out, channel11_Kernel53_Valid_Out, channel12_Kernel53_Valid_Out, channel13_Kernel53_Valid_Out, channel14_Kernel53_Valid_Out, channel15_Kernel53_Valid_Out, channel16_Kernel53_Valid_Out, channel17_Kernel53_Valid_Out, channel18_Kernel53_Valid_Out, channel19_Kernel53_Valid_Out, channel20_Kernel53_Valid_Out, channel21_Kernel53_Valid_Out, channel22_Kernel53_Valid_Out, channel23_Kernel53_Valid_Out, channel24_Kernel53_Valid_Out, channel25_Kernel53_Valid_Out, channel26_Kernel53_Valid_Out, channel27_Kernel53_Valid_Out, channel28_Kernel53_Valid_Out, channel29_Kernel53_Valid_Out, channel30_Kernel53_Valid_Out, channel31_Kernel53_Valid_Out, channel32_Kernel53_Valid_Out, channel33_Kernel53_Valid_Out, channel34_Kernel53_Valid_Out, channel35_Kernel53_Valid_Out, channel36_Kernel53_Valid_Out, channel37_Kernel53_Valid_Out, channel38_Kernel53_Valid_Out, channel39_Kernel53_Valid_Out, channel40_Kernel53_Valid_Out, channel41_Kernel53_Valid_Out, channel42_Kernel53_Valid_Out, channel43_Kernel53_Valid_Out, channel44_Kernel53_Valid_Out, channel45_Kernel53_Valid_Out, channel46_Kernel53_Valid_Out, channel47_Kernel53_Valid_Out, channel48_Kernel53_Valid_Out, channel49_Kernel53_Valid_Out, channel50_Kernel53_Valid_Out, channel51_Kernel53_Valid_Out, channel52_Kernel53_Valid_Out, channel53_Kernel53_Valid_Out, channel54_Kernel53_Valid_Out, channel55_Kernel53_Valid_Out, channel56_Kernel53_Valid_Out, channel57_Kernel53_Valid_Out, channel58_Kernel53_Valid_Out, channel59_Kernel53_Valid_Out, channel60_Kernel53_Valid_Out, channel61_Kernel53_Valid_Out, channel62_Kernel53_Valid_Out, channel63_Kernel53_Valid_Out, channel64_Kernel53_Valid_Out;

	assign add_kernel53=channel1_Kernel53_Valid_Out & channel2_Kernel53_Valid_Out & channel3_Kernel53_Valid_Out & channel4_Kernel53_Valid_Out & channel5_Kernel53_Valid_Out & channel6_Kernel53_Valid_Out & channel7_Kernel53_Valid_Out & channel8_Kernel53_Valid_Out & channel9_Kernel53_Valid_Out & channel10_Kernel53_Valid_Out & channel11_Kernel53_Valid_Out & channel12_Kernel53_Valid_Out & channel13_Kernel53_Valid_Out & channel14_Kernel53_Valid_Out & channel15_Kernel53_Valid_Out & channel16_Kernel53_Valid_Out & channel17_Kernel53_Valid_Out & channel18_Kernel53_Valid_Out & channel19_Kernel53_Valid_Out & channel20_Kernel53_Valid_Out & channel21_Kernel53_Valid_Out & channel22_Kernel53_Valid_Out & channel23_Kernel53_Valid_Out & channel24_Kernel53_Valid_Out & channel25_Kernel53_Valid_Out & channel26_Kernel53_Valid_Out & channel27_Kernel53_Valid_Out & channel28_Kernel53_Valid_Out & channel29_Kernel53_Valid_Out & channel30_Kernel53_Valid_Out & channel31_Kernel53_Valid_Out & channel32_Kernel53_Valid_Out & channel33_Kernel53_Valid_Out & channel34_Kernel53_Valid_Out & channel35_Kernel53_Valid_Out & channel36_Kernel53_Valid_Out & channel37_Kernel53_Valid_Out & channel38_Kernel53_Valid_Out & channel39_Kernel53_Valid_Out & channel40_Kernel53_Valid_Out & channel41_Kernel53_Valid_Out & channel42_Kernel53_Valid_Out & channel43_Kernel53_Valid_Out & channel44_Kernel53_Valid_Out & channel45_Kernel53_Valid_Out & channel46_Kernel53_Valid_Out & channel47_Kernel53_Valid_Out & channel48_Kernel53_Valid_Out & channel49_Kernel53_Valid_Out & channel50_Kernel53_Valid_Out & channel51_Kernel53_Valid_Out & channel52_Kernel53_Valid_Out & channel53_Kernel53_Valid_Out & channel54_Kernel53_Valid_Out & channel55_Kernel53_Valid_Out & channel56_Kernel53_Valid_Out & channel57_Kernel53_Valid_Out & channel58_Kernel53_Valid_Out & channel59_Kernel53_Valid_Out & channel60_Kernel53_Valid_Out & channel61_Kernel53_Valid_Out & channel62_Kernel53_Valid_Out & channel63_Kernel53_Valid_Out & channel64_Kernel53_Valid_Out;

	wire channel1_Kernel54_Valid_Out, channel2_Kernel54_Valid_Out, channel3_Kernel54_Valid_Out, channel4_Kernel54_Valid_Out, channel5_Kernel54_Valid_Out, channel6_Kernel54_Valid_Out, channel7_Kernel54_Valid_Out, channel8_Kernel54_Valid_Out, channel9_Kernel54_Valid_Out, channel10_Kernel54_Valid_Out, channel11_Kernel54_Valid_Out, channel12_Kernel54_Valid_Out, channel13_Kernel54_Valid_Out, channel14_Kernel54_Valid_Out, channel15_Kernel54_Valid_Out, channel16_Kernel54_Valid_Out, channel17_Kernel54_Valid_Out, channel18_Kernel54_Valid_Out, channel19_Kernel54_Valid_Out, channel20_Kernel54_Valid_Out, channel21_Kernel54_Valid_Out, channel22_Kernel54_Valid_Out, channel23_Kernel54_Valid_Out, channel24_Kernel54_Valid_Out, channel25_Kernel54_Valid_Out, channel26_Kernel54_Valid_Out, channel27_Kernel54_Valid_Out, channel28_Kernel54_Valid_Out, channel29_Kernel54_Valid_Out, channel30_Kernel54_Valid_Out, channel31_Kernel54_Valid_Out, channel32_Kernel54_Valid_Out, channel33_Kernel54_Valid_Out, channel34_Kernel54_Valid_Out, channel35_Kernel54_Valid_Out, channel36_Kernel54_Valid_Out, channel37_Kernel54_Valid_Out, channel38_Kernel54_Valid_Out, channel39_Kernel54_Valid_Out, channel40_Kernel54_Valid_Out, channel41_Kernel54_Valid_Out, channel42_Kernel54_Valid_Out, channel43_Kernel54_Valid_Out, channel44_Kernel54_Valid_Out, channel45_Kernel54_Valid_Out, channel46_Kernel54_Valid_Out, channel47_Kernel54_Valid_Out, channel48_Kernel54_Valid_Out, channel49_Kernel54_Valid_Out, channel50_Kernel54_Valid_Out, channel51_Kernel54_Valid_Out, channel52_Kernel54_Valid_Out, channel53_Kernel54_Valid_Out, channel54_Kernel54_Valid_Out, channel55_Kernel54_Valid_Out, channel56_Kernel54_Valid_Out, channel57_Kernel54_Valid_Out, channel58_Kernel54_Valid_Out, channel59_Kernel54_Valid_Out, channel60_Kernel54_Valid_Out, channel61_Kernel54_Valid_Out, channel62_Kernel54_Valid_Out, channel63_Kernel54_Valid_Out, channel64_Kernel54_Valid_Out;

	assign add_kernel54=channel1_Kernel54_Valid_Out & channel2_Kernel54_Valid_Out & channel3_Kernel54_Valid_Out & channel4_Kernel54_Valid_Out & channel5_Kernel54_Valid_Out & channel6_Kernel54_Valid_Out & channel7_Kernel54_Valid_Out & channel8_Kernel54_Valid_Out & channel9_Kernel54_Valid_Out & channel10_Kernel54_Valid_Out & channel11_Kernel54_Valid_Out & channel12_Kernel54_Valid_Out & channel13_Kernel54_Valid_Out & channel14_Kernel54_Valid_Out & channel15_Kernel54_Valid_Out & channel16_Kernel54_Valid_Out & channel17_Kernel54_Valid_Out & channel18_Kernel54_Valid_Out & channel19_Kernel54_Valid_Out & channel20_Kernel54_Valid_Out & channel21_Kernel54_Valid_Out & channel22_Kernel54_Valid_Out & channel23_Kernel54_Valid_Out & channel24_Kernel54_Valid_Out & channel25_Kernel54_Valid_Out & channel26_Kernel54_Valid_Out & channel27_Kernel54_Valid_Out & channel28_Kernel54_Valid_Out & channel29_Kernel54_Valid_Out & channel30_Kernel54_Valid_Out & channel31_Kernel54_Valid_Out & channel32_Kernel54_Valid_Out & channel33_Kernel54_Valid_Out & channel34_Kernel54_Valid_Out & channel35_Kernel54_Valid_Out & channel36_Kernel54_Valid_Out & channel37_Kernel54_Valid_Out & channel38_Kernel54_Valid_Out & channel39_Kernel54_Valid_Out & channel40_Kernel54_Valid_Out & channel41_Kernel54_Valid_Out & channel42_Kernel54_Valid_Out & channel43_Kernel54_Valid_Out & channel44_Kernel54_Valid_Out & channel45_Kernel54_Valid_Out & channel46_Kernel54_Valid_Out & channel47_Kernel54_Valid_Out & channel48_Kernel54_Valid_Out & channel49_Kernel54_Valid_Out & channel50_Kernel54_Valid_Out & channel51_Kernel54_Valid_Out & channel52_Kernel54_Valid_Out & channel53_Kernel54_Valid_Out & channel54_Kernel54_Valid_Out & channel55_Kernel54_Valid_Out & channel56_Kernel54_Valid_Out & channel57_Kernel54_Valid_Out & channel58_Kernel54_Valid_Out & channel59_Kernel54_Valid_Out & channel60_Kernel54_Valid_Out & channel61_Kernel54_Valid_Out & channel62_Kernel54_Valid_Out & channel63_Kernel54_Valid_Out & channel64_Kernel54_Valid_Out;

	wire channel1_Kernel55_Valid_Out, channel2_Kernel55_Valid_Out, channel3_Kernel55_Valid_Out, channel4_Kernel55_Valid_Out, channel5_Kernel55_Valid_Out, channel6_Kernel55_Valid_Out, channel7_Kernel55_Valid_Out, channel8_Kernel55_Valid_Out, channel9_Kernel55_Valid_Out, channel10_Kernel55_Valid_Out, channel11_Kernel55_Valid_Out, channel12_Kernel55_Valid_Out, channel13_Kernel55_Valid_Out, channel14_Kernel55_Valid_Out, channel15_Kernel55_Valid_Out, channel16_Kernel55_Valid_Out, channel17_Kernel55_Valid_Out, channel18_Kernel55_Valid_Out, channel19_Kernel55_Valid_Out, channel20_Kernel55_Valid_Out, channel21_Kernel55_Valid_Out, channel22_Kernel55_Valid_Out, channel23_Kernel55_Valid_Out, channel24_Kernel55_Valid_Out, channel25_Kernel55_Valid_Out, channel26_Kernel55_Valid_Out, channel27_Kernel55_Valid_Out, channel28_Kernel55_Valid_Out, channel29_Kernel55_Valid_Out, channel30_Kernel55_Valid_Out, channel31_Kernel55_Valid_Out, channel32_Kernel55_Valid_Out, channel33_Kernel55_Valid_Out, channel34_Kernel55_Valid_Out, channel35_Kernel55_Valid_Out, channel36_Kernel55_Valid_Out, channel37_Kernel55_Valid_Out, channel38_Kernel55_Valid_Out, channel39_Kernel55_Valid_Out, channel40_Kernel55_Valid_Out, channel41_Kernel55_Valid_Out, channel42_Kernel55_Valid_Out, channel43_Kernel55_Valid_Out, channel44_Kernel55_Valid_Out, channel45_Kernel55_Valid_Out, channel46_Kernel55_Valid_Out, channel47_Kernel55_Valid_Out, channel48_Kernel55_Valid_Out, channel49_Kernel55_Valid_Out, channel50_Kernel55_Valid_Out, channel51_Kernel55_Valid_Out, channel52_Kernel55_Valid_Out, channel53_Kernel55_Valid_Out, channel54_Kernel55_Valid_Out, channel55_Kernel55_Valid_Out, channel56_Kernel55_Valid_Out, channel57_Kernel55_Valid_Out, channel58_Kernel55_Valid_Out, channel59_Kernel55_Valid_Out, channel60_Kernel55_Valid_Out, channel61_Kernel55_Valid_Out, channel62_Kernel55_Valid_Out, channel63_Kernel55_Valid_Out, channel64_Kernel55_Valid_Out;

	assign add_kernel55=channel1_Kernel55_Valid_Out & channel2_Kernel55_Valid_Out & channel3_Kernel55_Valid_Out & channel4_Kernel55_Valid_Out & channel5_Kernel55_Valid_Out & channel6_Kernel55_Valid_Out & channel7_Kernel55_Valid_Out & channel8_Kernel55_Valid_Out & channel9_Kernel55_Valid_Out & channel10_Kernel55_Valid_Out & channel11_Kernel55_Valid_Out & channel12_Kernel55_Valid_Out & channel13_Kernel55_Valid_Out & channel14_Kernel55_Valid_Out & channel15_Kernel55_Valid_Out & channel16_Kernel55_Valid_Out & channel17_Kernel55_Valid_Out & channel18_Kernel55_Valid_Out & channel19_Kernel55_Valid_Out & channel20_Kernel55_Valid_Out & channel21_Kernel55_Valid_Out & channel22_Kernel55_Valid_Out & channel23_Kernel55_Valid_Out & channel24_Kernel55_Valid_Out & channel25_Kernel55_Valid_Out & channel26_Kernel55_Valid_Out & channel27_Kernel55_Valid_Out & channel28_Kernel55_Valid_Out & channel29_Kernel55_Valid_Out & channel30_Kernel55_Valid_Out & channel31_Kernel55_Valid_Out & channel32_Kernel55_Valid_Out & channel33_Kernel55_Valid_Out & channel34_Kernel55_Valid_Out & channel35_Kernel55_Valid_Out & channel36_Kernel55_Valid_Out & channel37_Kernel55_Valid_Out & channel38_Kernel55_Valid_Out & channel39_Kernel55_Valid_Out & channel40_Kernel55_Valid_Out & channel41_Kernel55_Valid_Out & channel42_Kernel55_Valid_Out & channel43_Kernel55_Valid_Out & channel44_Kernel55_Valid_Out & channel45_Kernel55_Valid_Out & channel46_Kernel55_Valid_Out & channel47_Kernel55_Valid_Out & channel48_Kernel55_Valid_Out & channel49_Kernel55_Valid_Out & channel50_Kernel55_Valid_Out & channel51_Kernel55_Valid_Out & channel52_Kernel55_Valid_Out & channel53_Kernel55_Valid_Out & channel54_Kernel55_Valid_Out & channel55_Kernel55_Valid_Out & channel56_Kernel55_Valid_Out & channel57_Kernel55_Valid_Out & channel58_Kernel55_Valid_Out & channel59_Kernel55_Valid_Out & channel60_Kernel55_Valid_Out & channel61_Kernel55_Valid_Out & channel62_Kernel55_Valid_Out & channel63_Kernel55_Valid_Out & channel64_Kernel55_Valid_Out;

	wire channel1_Kernel56_Valid_Out, channel2_Kernel56_Valid_Out, channel3_Kernel56_Valid_Out, channel4_Kernel56_Valid_Out, channel5_Kernel56_Valid_Out, channel6_Kernel56_Valid_Out, channel7_Kernel56_Valid_Out, channel8_Kernel56_Valid_Out, channel9_Kernel56_Valid_Out, channel10_Kernel56_Valid_Out, channel11_Kernel56_Valid_Out, channel12_Kernel56_Valid_Out, channel13_Kernel56_Valid_Out, channel14_Kernel56_Valid_Out, channel15_Kernel56_Valid_Out, channel16_Kernel56_Valid_Out, channel17_Kernel56_Valid_Out, channel18_Kernel56_Valid_Out, channel19_Kernel56_Valid_Out, channel20_Kernel56_Valid_Out, channel21_Kernel56_Valid_Out, channel22_Kernel56_Valid_Out, channel23_Kernel56_Valid_Out, channel24_Kernel56_Valid_Out, channel25_Kernel56_Valid_Out, channel26_Kernel56_Valid_Out, channel27_Kernel56_Valid_Out, channel28_Kernel56_Valid_Out, channel29_Kernel56_Valid_Out, channel30_Kernel56_Valid_Out, channel31_Kernel56_Valid_Out, channel32_Kernel56_Valid_Out, channel33_Kernel56_Valid_Out, channel34_Kernel56_Valid_Out, channel35_Kernel56_Valid_Out, channel36_Kernel56_Valid_Out, channel37_Kernel56_Valid_Out, channel38_Kernel56_Valid_Out, channel39_Kernel56_Valid_Out, channel40_Kernel56_Valid_Out, channel41_Kernel56_Valid_Out, channel42_Kernel56_Valid_Out, channel43_Kernel56_Valid_Out, channel44_Kernel56_Valid_Out, channel45_Kernel56_Valid_Out, channel46_Kernel56_Valid_Out, channel47_Kernel56_Valid_Out, channel48_Kernel56_Valid_Out, channel49_Kernel56_Valid_Out, channel50_Kernel56_Valid_Out, channel51_Kernel56_Valid_Out, channel52_Kernel56_Valid_Out, channel53_Kernel56_Valid_Out, channel54_Kernel56_Valid_Out, channel55_Kernel56_Valid_Out, channel56_Kernel56_Valid_Out, channel57_Kernel56_Valid_Out, channel58_Kernel56_Valid_Out, channel59_Kernel56_Valid_Out, channel60_Kernel56_Valid_Out, channel61_Kernel56_Valid_Out, channel62_Kernel56_Valid_Out, channel63_Kernel56_Valid_Out, channel64_Kernel56_Valid_Out;

	assign add_kernel56=channel1_Kernel56_Valid_Out & channel2_Kernel56_Valid_Out & channel3_Kernel56_Valid_Out & channel4_Kernel56_Valid_Out & channel5_Kernel56_Valid_Out & channel6_Kernel56_Valid_Out & channel7_Kernel56_Valid_Out & channel8_Kernel56_Valid_Out & channel9_Kernel56_Valid_Out & channel10_Kernel56_Valid_Out & channel11_Kernel56_Valid_Out & channel12_Kernel56_Valid_Out & channel13_Kernel56_Valid_Out & channel14_Kernel56_Valid_Out & channel15_Kernel56_Valid_Out & channel16_Kernel56_Valid_Out & channel17_Kernel56_Valid_Out & channel18_Kernel56_Valid_Out & channel19_Kernel56_Valid_Out & channel20_Kernel56_Valid_Out & channel21_Kernel56_Valid_Out & channel22_Kernel56_Valid_Out & channel23_Kernel56_Valid_Out & channel24_Kernel56_Valid_Out & channel25_Kernel56_Valid_Out & channel26_Kernel56_Valid_Out & channel27_Kernel56_Valid_Out & channel28_Kernel56_Valid_Out & channel29_Kernel56_Valid_Out & channel30_Kernel56_Valid_Out & channel31_Kernel56_Valid_Out & channel32_Kernel56_Valid_Out & channel33_Kernel56_Valid_Out & channel34_Kernel56_Valid_Out & channel35_Kernel56_Valid_Out & channel36_Kernel56_Valid_Out & channel37_Kernel56_Valid_Out & channel38_Kernel56_Valid_Out & channel39_Kernel56_Valid_Out & channel40_Kernel56_Valid_Out & channel41_Kernel56_Valid_Out & channel42_Kernel56_Valid_Out & channel43_Kernel56_Valid_Out & channel44_Kernel56_Valid_Out & channel45_Kernel56_Valid_Out & channel46_Kernel56_Valid_Out & channel47_Kernel56_Valid_Out & channel48_Kernel56_Valid_Out & channel49_Kernel56_Valid_Out & channel50_Kernel56_Valid_Out & channel51_Kernel56_Valid_Out & channel52_Kernel56_Valid_Out & channel53_Kernel56_Valid_Out & channel54_Kernel56_Valid_Out & channel55_Kernel56_Valid_Out & channel56_Kernel56_Valid_Out & channel57_Kernel56_Valid_Out & channel58_Kernel56_Valid_Out & channel59_Kernel56_Valid_Out & channel60_Kernel56_Valid_Out & channel61_Kernel56_Valid_Out & channel62_Kernel56_Valid_Out & channel63_Kernel56_Valid_Out & channel64_Kernel56_Valid_Out;

	wire channel1_Kernel57_Valid_Out, channel2_Kernel57_Valid_Out, channel3_Kernel57_Valid_Out, channel4_Kernel57_Valid_Out, channel5_Kernel57_Valid_Out, channel6_Kernel57_Valid_Out, channel7_Kernel57_Valid_Out, channel8_Kernel57_Valid_Out, channel9_Kernel57_Valid_Out, channel10_Kernel57_Valid_Out, channel11_Kernel57_Valid_Out, channel12_Kernel57_Valid_Out, channel13_Kernel57_Valid_Out, channel14_Kernel57_Valid_Out, channel15_Kernel57_Valid_Out, channel16_Kernel57_Valid_Out, channel17_Kernel57_Valid_Out, channel18_Kernel57_Valid_Out, channel19_Kernel57_Valid_Out, channel20_Kernel57_Valid_Out, channel21_Kernel57_Valid_Out, channel22_Kernel57_Valid_Out, channel23_Kernel57_Valid_Out, channel24_Kernel57_Valid_Out, channel25_Kernel57_Valid_Out, channel26_Kernel57_Valid_Out, channel27_Kernel57_Valid_Out, channel28_Kernel57_Valid_Out, channel29_Kernel57_Valid_Out, channel30_Kernel57_Valid_Out, channel31_Kernel57_Valid_Out, channel32_Kernel57_Valid_Out, channel33_Kernel57_Valid_Out, channel34_Kernel57_Valid_Out, channel35_Kernel57_Valid_Out, channel36_Kernel57_Valid_Out, channel37_Kernel57_Valid_Out, channel38_Kernel57_Valid_Out, channel39_Kernel57_Valid_Out, channel40_Kernel57_Valid_Out, channel41_Kernel57_Valid_Out, channel42_Kernel57_Valid_Out, channel43_Kernel57_Valid_Out, channel44_Kernel57_Valid_Out, channel45_Kernel57_Valid_Out, channel46_Kernel57_Valid_Out, channel47_Kernel57_Valid_Out, channel48_Kernel57_Valid_Out, channel49_Kernel57_Valid_Out, channel50_Kernel57_Valid_Out, channel51_Kernel57_Valid_Out, channel52_Kernel57_Valid_Out, channel53_Kernel57_Valid_Out, channel54_Kernel57_Valid_Out, channel55_Kernel57_Valid_Out, channel56_Kernel57_Valid_Out, channel57_Kernel57_Valid_Out, channel58_Kernel57_Valid_Out, channel59_Kernel57_Valid_Out, channel60_Kernel57_Valid_Out, channel61_Kernel57_Valid_Out, channel62_Kernel57_Valid_Out, channel63_Kernel57_Valid_Out, channel64_Kernel57_Valid_Out;

	assign add_kernel57=channel1_Kernel57_Valid_Out & channel2_Kernel57_Valid_Out & channel3_Kernel57_Valid_Out & channel4_Kernel57_Valid_Out & channel5_Kernel57_Valid_Out & channel6_Kernel57_Valid_Out & channel7_Kernel57_Valid_Out & channel8_Kernel57_Valid_Out & channel9_Kernel57_Valid_Out & channel10_Kernel57_Valid_Out & channel11_Kernel57_Valid_Out & channel12_Kernel57_Valid_Out & channel13_Kernel57_Valid_Out & channel14_Kernel57_Valid_Out & channel15_Kernel57_Valid_Out & channel16_Kernel57_Valid_Out & channel17_Kernel57_Valid_Out & channel18_Kernel57_Valid_Out & channel19_Kernel57_Valid_Out & channel20_Kernel57_Valid_Out & channel21_Kernel57_Valid_Out & channel22_Kernel57_Valid_Out & channel23_Kernel57_Valid_Out & channel24_Kernel57_Valid_Out & channel25_Kernel57_Valid_Out & channel26_Kernel57_Valid_Out & channel27_Kernel57_Valid_Out & channel28_Kernel57_Valid_Out & channel29_Kernel57_Valid_Out & channel30_Kernel57_Valid_Out & channel31_Kernel57_Valid_Out & channel32_Kernel57_Valid_Out & channel33_Kernel57_Valid_Out & channel34_Kernel57_Valid_Out & channel35_Kernel57_Valid_Out & channel36_Kernel57_Valid_Out & channel37_Kernel57_Valid_Out & channel38_Kernel57_Valid_Out & channel39_Kernel57_Valid_Out & channel40_Kernel57_Valid_Out & channel41_Kernel57_Valid_Out & channel42_Kernel57_Valid_Out & channel43_Kernel57_Valid_Out & channel44_Kernel57_Valid_Out & channel45_Kernel57_Valid_Out & channel46_Kernel57_Valid_Out & channel47_Kernel57_Valid_Out & channel48_Kernel57_Valid_Out & channel49_Kernel57_Valid_Out & channel50_Kernel57_Valid_Out & channel51_Kernel57_Valid_Out & channel52_Kernel57_Valid_Out & channel53_Kernel57_Valid_Out & channel54_Kernel57_Valid_Out & channel55_Kernel57_Valid_Out & channel56_Kernel57_Valid_Out & channel57_Kernel57_Valid_Out & channel58_Kernel57_Valid_Out & channel59_Kernel57_Valid_Out & channel60_Kernel57_Valid_Out & channel61_Kernel57_Valid_Out & channel62_Kernel57_Valid_Out & channel63_Kernel57_Valid_Out & channel64_Kernel57_Valid_Out;

	wire channel1_Kernel58_Valid_Out, channel2_Kernel58_Valid_Out, channel3_Kernel58_Valid_Out, channel4_Kernel58_Valid_Out, channel5_Kernel58_Valid_Out, channel6_Kernel58_Valid_Out, channel7_Kernel58_Valid_Out, channel8_Kernel58_Valid_Out, channel9_Kernel58_Valid_Out, channel10_Kernel58_Valid_Out, channel11_Kernel58_Valid_Out, channel12_Kernel58_Valid_Out, channel13_Kernel58_Valid_Out, channel14_Kernel58_Valid_Out, channel15_Kernel58_Valid_Out, channel16_Kernel58_Valid_Out, channel17_Kernel58_Valid_Out, channel18_Kernel58_Valid_Out, channel19_Kernel58_Valid_Out, channel20_Kernel58_Valid_Out, channel21_Kernel58_Valid_Out, channel22_Kernel58_Valid_Out, channel23_Kernel58_Valid_Out, channel24_Kernel58_Valid_Out, channel25_Kernel58_Valid_Out, channel26_Kernel58_Valid_Out, channel27_Kernel58_Valid_Out, channel28_Kernel58_Valid_Out, channel29_Kernel58_Valid_Out, channel30_Kernel58_Valid_Out, channel31_Kernel58_Valid_Out, channel32_Kernel58_Valid_Out, channel33_Kernel58_Valid_Out, channel34_Kernel58_Valid_Out, channel35_Kernel58_Valid_Out, channel36_Kernel58_Valid_Out, channel37_Kernel58_Valid_Out, channel38_Kernel58_Valid_Out, channel39_Kernel58_Valid_Out, channel40_Kernel58_Valid_Out, channel41_Kernel58_Valid_Out, channel42_Kernel58_Valid_Out, channel43_Kernel58_Valid_Out, channel44_Kernel58_Valid_Out, channel45_Kernel58_Valid_Out, channel46_Kernel58_Valid_Out, channel47_Kernel58_Valid_Out, channel48_Kernel58_Valid_Out, channel49_Kernel58_Valid_Out, channel50_Kernel58_Valid_Out, channel51_Kernel58_Valid_Out, channel52_Kernel58_Valid_Out, channel53_Kernel58_Valid_Out, channel54_Kernel58_Valid_Out, channel55_Kernel58_Valid_Out, channel56_Kernel58_Valid_Out, channel57_Kernel58_Valid_Out, channel58_Kernel58_Valid_Out, channel59_Kernel58_Valid_Out, channel60_Kernel58_Valid_Out, channel61_Kernel58_Valid_Out, channel62_Kernel58_Valid_Out, channel63_Kernel58_Valid_Out, channel64_Kernel58_Valid_Out;

	assign add_kernel58=channel1_Kernel58_Valid_Out & channel2_Kernel58_Valid_Out & channel3_Kernel58_Valid_Out & channel4_Kernel58_Valid_Out & channel5_Kernel58_Valid_Out & channel6_Kernel58_Valid_Out & channel7_Kernel58_Valid_Out & channel8_Kernel58_Valid_Out & channel9_Kernel58_Valid_Out & channel10_Kernel58_Valid_Out & channel11_Kernel58_Valid_Out & channel12_Kernel58_Valid_Out & channel13_Kernel58_Valid_Out & channel14_Kernel58_Valid_Out & channel15_Kernel58_Valid_Out & channel16_Kernel58_Valid_Out & channel17_Kernel58_Valid_Out & channel18_Kernel58_Valid_Out & channel19_Kernel58_Valid_Out & channel20_Kernel58_Valid_Out & channel21_Kernel58_Valid_Out & channel22_Kernel58_Valid_Out & channel23_Kernel58_Valid_Out & channel24_Kernel58_Valid_Out & channel25_Kernel58_Valid_Out & channel26_Kernel58_Valid_Out & channel27_Kernel58_Valid_Out & channel28_Kernel58_Valid_Out & channel29_Kernel58_Valid_Out & channel30_Kernel58_Valid_Out & channel31_Kernel58_Valid_Out & channel32_Kernel58_Valid_Out & channel33_Kernel58_Valid_Out & channel34_Kernel58_Valid_Out & channel35_Kernel58_Valid_Out & channel36_Kernel58_Valid_Out & channel37_Kernel58_Valid_Out & channel38_Kernel58_Valid_Out & channel39_Kernel58_Valid_Out & channel40_Kernel58_Valid_Out & channel41_Kernel58_Valid_Out & channel42_Kernel58_Valid_Out & channel43_Kernel58_Valid_Out & channel44_Kernel58_Valid_Out & channel45_Kernel58_Valid_Out & channel46_Kernel58_Valid_Out & channel47_Kernel58_Valid_Out & channel48_Kernel58_Valid_Out & channel49_Kernel58_Valid_Out & channel50_Kernel58_Valid_Out & channel51_Kernel58_Valid_Out & channel52_Kernel58_Valid_Out & channel53_Kernel58_Valid_Out & channel54_Kernel58_Valid_Out & channel55_Kernel58_Valid_Out & channel56_Kernel58_Valid_Out & channel57_Kernel58_Valid_Out & channel58_Kernel58_Valid_Out & channel59_Kernel58_Valid_Out & channel60_Kernel58_Valid_Out & channel61_Kernel58_Valid_Out & channel62_Kernel58_Valid_Out & channel63_Kernel58_Valid_Out & channel64_Kernel58_Valid_Out;

	wire channel1_Kernel59_Valid_Out, channel2_Kernel59_Valid_Out, channel3_Kernel59_Valid_Out, channel4_Kernel59_Valid_Out, channel5_Kernel59_Valid_Out, channel6_Kernel59_Valid_Out, channel7_Kernel59_Valid_Out, channel8_Kernel59_Valid_Out, channel9_Kernel59_Valid_Out, channel10_Kernel59_Valid_Out, channel11_Kernel59_Valid_Out, channel12_Kernel59_Valid_Out, channel13_Kernel59_Valid_Out, channel14_Kernel59_Valid_Out, channel15_Kernel59_Valid_Out, channel16_Kernel59_Valid_Out, channel17_Kernel59_Valid_Out, channel18_Kernel59_Valid_Out, channel19_Kernel59_Valid_Out, channel20_Kernel59_Valid_Out, channel21_Kernel59_Valid_Out, channel22_Kernel59_Valid_Out, channel23_Kernel59_Valid_Out, channel24_Kernel59_Valid_Out, channel25_Kernel59_Valid_Out, channel26_Kernel59_Valid_Out, channel27_Kernel59_Valid_Out, channel28_Kernel59_Valid_Out, channel29_Kernel59_Valid_Out, channel30_Kernel59_Valid_Out, channel31_Kernel59_Valid_Out, channel32_Kernel59_Valid_Out, channel33_Kernel59_Valid_Out, channel34_Kernel59_Valid_Out, channel35_Kernel59_Valid_Out, channel36_Kernel59_Valid_Out, channel37_Kernel59_Valid_Out, channel38_Kernel59_Valid_Out, channel39_Kernel59_Valid_Out, channel40_Kernel59_Valid_Out, channel41_Kernel59_Valid_Out, channel42_Kernel59_Valid_Out, channel43_Kernel59_Valid_Out, channel44_Kernel59_Valid_Out, channel45_Kernel59_Valid_Out, channel46_Kernel59_Valid_Out, channel47_Kernel59_Valid_Out, channel48_Kernel59_Valid_Out, channel49_Kernel59_Valid_Out, channel50_Kernel59_Valid_Out, channel51_Kernel59_Valid_Out, channel52_Kernel59_Valid_Out, channel53_Kernel59_Valid_Out, channel54_Kernel59_Valid_Out, channel55_Kernel59_Valid_Out, channel56_Kernel59_Valid_Out, channel57_Kernel59_Valid_Out, channel58_Kernel59_Valid_Out, channel59_Kernel59_Valid_Out, channel60_Kernel59_Valid_Out, channel61_Kernel59_Valid_Out, channel62_Kernel59_Valid_Out, channel63_Kernel59_Valid_Out, channel64_Kernel59_Valid_Out;

	assign add_kernel59=channel1_Kernel59_Valid_Out & channel2_Kernel59_Valid_Out & channel3_Kernel59_Valid_Out & channel4_Kernel59_Valid_Out & channel5_Kernel59_Valid_Out & channel6_Kernel59_Valid_Out & channel7_Kernel59_Valid_Out & channel8_Kernel59_Valid_Out & channel9_Kernel59_Valid_Out & channel10_Kernel59_Valid_Out & channel11_Kernel59_Valid_Out & channel12_Kernel59_Valid_Out & channel13_Kernel59_Valid_Out & channel14_Kernel59_Valid_Out & channel15_Kernel59_Valid_Out & channel16_Kernel59_Valid_Out & channel17_Kernel59_Valid_Out & channel18_Kernel59_Valid_Out & channel19_Kernel59_Valid_Out & channel20_Kernel59_Valid_Out & channel21_Kernel59_Valid_Out & channel22_Kernel59_Valid_Out & channel23_Kernel59_Valid_Out & channel24_Kernel59_Valid_Out & channel25_Kernel59_Valid_Out & channel26_Kernel59_Valid_Out & channel27_Kernel59_Valid_Out & channel28_Kernel59_Valid_Out & channel29_Kernel59_Valid_Out & channel30_Kernel59_Valid_Out & channel31_Kernel59_Valid_Out & channel32_Kernel59_Valid_Out & channel33_Kernel59_Valid_Out & channel34_Kernel59_Valid_Out & channel35_Kernel59_Valid_Out & channel36_Kernel59_Valid_Out & channel37_Kernel59_Valid_Out & channel38_Kernel59_Valid_Out & channel39_Kernel59_Valid_Out & channel40_Kernel59_Valid_Out & channel41_Kernel59_Valid_Out & channel42_Kernel59_Valid_Out & channel43_Kernel59_Valid_Out & channel44_Kernel59_Valid_Out & channel45_Kernel59_Valid_Out & channel46_Kernel59_Valid_Out & channel47_Kernel59_Valid_Out & channel48_Kernel59_Valid_Out & channel49_Kernel59_Valid_Out & channel50_Kernel59_Valid_Out & channel51_Kernel59_Valid_Out & channel52_Kernel59_Valid_Out & channel53_Kernel59_Valid_Out & channel54_Kernel59_Valid_Out & channel55_Kernel59_Valid_Out & channel56_Kernel59_Valid_Out & channel57_Kernel59_Valid_Out & channel58_Kernel59_Valid_Out & channel59_Kernel59_Valid_Out & channel60_Kernel59_Valid_Out & channel61_Kernel59_Valid_Out & channel62_Kernel59_Valid_Out & channel63_Kernel59_Valid_Out & channel64_Kernel59_Valid_Out;

	wire channel1_Kernel60_Valid_Out, channel2_Kernel60_Valid_Out, channel3_Kernel60_Valid_Out, channel4_Kernel60_Valid_Out, channel5_Kernel60_Valid_Out, channel6_Kernel60_Valid_Out, channel7_Kernel60_Valid_Out, channel8_Kernel60_Valid_Out, channel9_Kernel60_Valid_Out, channel10_Kernel60_Valid_Out, channel11_Kernel60_Valid_Out, channel12_Kernel60_Valid_Out, channel13_Kernel60_Valid_Out, channel14_Kernel60_Valid_Out, channel15_Kernel60_Valid_Out, channel16_Kernel60_Valid_Out, channel17_Kernel60_Valid_Out, channel18_Kernel60_Valid_Out, channel19_Kernel60_Valid_Out, channel20_Kernel60_Valid_Out, channel21_Kernel60_Valid_Out, channel22_Kernel60_Valid_Out, channel23_Kernel60_Valid_Out, channel24_Kernel60_Valid_Out, channel25_Kernel60_Valid_Out, channel26_Kernel60_Valid_Out, channel27_Kernel60_Valid_Out, channel28_Kernel60_Valid_Out, channel29_Kernel60_Valid_Out, channel30_Kernel60_Valid_Out, channel31_Kernel60_Valid_Out, channel32_Kernel60_Valid_Out, channel33_Kernel60_Valid_Out, channel34_Kernel60_Valid_Out, channel35_Kernel60_Valid_Out, channel36_Kernel60_Valid_Out, channel37_Kernel60_Valid_Out, channel38_Kernel60_Valid_Out, channel39_Kernel60_Valid_Out, channel40_Kernel60_Valid_Out, channel41_Kernel60_Valid_Out, channel42_Kernel60_Valid_Out, channel43_Kernel60_Valid_Out, channel44_Kernel60_Valid_Out, channel45_Kernel60_Valid_Out, channel46_Kernel60_Valid_Out, channel47_Kernel60_Valid_Out, channel48_Kernel60_Valid_Out, channel49_Kernel60_Valid_Out, channel50_Kernel60_Valid_Out, channel51_Kernel60_Valid_Out, channel52_Kernel60_Valid_Out, channel53_Kernel60_Valid_Out, channel54_Kernel60_Valid_Out, channel55_Kernel60_Valid_Out, channel56_Kernel60_Valid_Out, channel57_Kernel60_Valid_Out, channel58_Kernel60_Valid_Out, channel59_Kernel60_Valid_Out, channel60_Kernel60_Valid_Out, channel61_Kernel60_Valid_Out, channel62_Kernel60_Valid_Out, channel63_Kernel60_Valid_Out, channel64_Kernel60_Valid_Out;

	assign add_kernel60=channel1_Kernel60_Valid_Out & channel2_Kernel60_Valid_Out & channel3_Kernel60_Valid_Out & channel4_Kernel60_Valid_Out & channel5_Kernel60_Valid_Out & channel6_Kernel60_Valid_Out & channel7_Kernel60_Valid_Out & channel8_Kernel60_Valid_Out & channel9_Kernel60_Valid_Out & channel10_Kernel60_Valid_Out & channel11_Kernel60_Valid_Out & channel12_Kernel60_Valid_Out & channel13_Kernel60_Valid_Out & channel14_Kernel60_Valid_Out & channel15_Kernel60_Valid_Out & channel16_Kernel60_Valid_Out & channel17_Kernel60_Valid_Out & channel18_Kernel60_Valid_Out & channel19_Kernel60_Valid_Out & channel20_Kernel60_Valid_Out & channel21_Kernel60_Valid_Out & channel22_Kernel60_Valid_Out & channel23_Kernel60_Valid_Out & channel24_Kernel60_Valid_Out & channel25_Kernel60_Valid_Out & channel26_Kernel60_Valid_Out & channel27_Kernel60_Valid_Out & channel28_Kernel60_Valid_Out & channel29_Kernel60_Valid_Out & channel30_Kernel60_Valid_Out & channel31_Kernel60_Valid_Out & channel32_Kernel60_Valid_Out & channel33_Kernel60_Valid_Out & channel34_Kernel60_Valid_Out & channel35_Kernel60_Valid_Out & channel36_Kernel60_Valid_Out & channel37_Kernel60_Valid_Out & channel38_Kernel60_Valid_Out & channel39_Kernel60_Valid_Out & channel40_Kernel60_Valid_Out & channel41_Kernel60_Valid_Out & channel42_Kernel60_Valid_Out & channel43_Kernel60_Valid_Out & channel44_Kernel60_Valid_Out & channel45_Kernel60_Valid_Out & channel46_Kernel60_Valid_Out & channel47_Kernel60_Valid_Out & channel48_Kernel60_Valid_Out & channel49_Kernel60_Valid_Out & channel50_Kernel60_Valid_Out & channel51_Kernel60_Valid_Out & channel52_Kernel60_Valid_Out & channel53_Kernel60_Valid_Out & channel54_Kernel60_Valid_Out & channel55_Kernel60_Valid_Out & channel56_Kernel60_Valid_Out & channel57_Kernel60_Valid_Out & channel58_Kernel60_Valid_Out & channel59_Kernel60_Valid_Out & channel60_Kernel60_Valid_Out & channel61_Kernel60_Valid_Out & channel62_Kernel60_Valid_Out & channel63_Kernel60_Valid_Out & channel64_Kernel60_Valid_Out;

	wire channel1_Kernel61_Valid_Out, channel2_Kernel61_Valid_Out, channel3_Kernel61_Valid_Out, channel4_Kernel61_Valid_Out, channel5_Kernel61_Valid_Out, channel6_Kernel61_Valid_Out, channel7_Kernel61_Valid_Out, channel8_Kernel61_Valid_Out, channel9_Kernel61_Valid_Out, channel10_Kernel61_Valid_Out, channel11_Kernel61_Valid_Out, channel12_Kernel61_Valid_Out, channel13_Kernel61_Valid_Out, channel14_Kernel61_Valid_Out, channel15_Kernel61_Valid_Out, channel16_Kernel61_Valid_Out, channel17_Kernel61_Valid_Out, channel18_Kernel61_Valid_Out, channel19_Kernel61_Valid_Out, channel20_Kernel61_Valid_Out, channel21_Kernel61_Valid_Out, channel22_Kernel61_Valid_Out, channel23_Kernel61_Valid_Out, channel24_Kernel61_Valid_Out, channel25_Kernel61_Valid_Out, channel26_Kernel61_Valid_Out, channel27_Kernel61_Valid_Out, channel28_Kernel61_Valid_Out, channel29_Kernel61_Valid_Out, channel30_Kernel61_Valid_Out, channel31_Kernel61_Valid_Out, channel32_Kernel61_Valid_Out, channel33_Kernel61_Valid_Out, channel34_Kernel61_Valid_Out, channel35_Kernel61_Valid_Out, channel36_Kernel61_Valid_Out, channel37_Kernel61_Valid_Out, channel38_Kernel61_Valid_Out, channel39_Kernel61_Valid_Out, channel40_Kernel61_Valid_Out, channel41_Kernel61_Valid_Out, channel42_Kernel61_Valid_Out, channel43_Kernel61_Valid_Out, channel44_Kernel61_Valid_Out, channel45_Kernel61_Valid_Out, channel46_Kernel61_Valid_Out, channel47_Kernel61_Valid_Out, channel48_Kernel61_Valid_Out, channel49_Kernel61_Valid_Out, channel50_Kernel61_Valid_Out, channel51_Kernel61_Valid_Out, channel52_Kernel61_Valid_Out, channel53_Kernel61_Valid_Out, channel54_Kernel61_Valid_Out, channel55_Kernel61_Valid_Out, channel56_Kernel61_Valid_Out, channel57_Kernel61_Valid_Out, channel58_Kernel61_Valid_Out, channel59_Kernel61_Valid_Out, channel60_Kernel61_Valid_Out, channel61_Kernel61_Valid_Out, channel62_Kernel61_Valid_Out, channel63_Kernel61_Valid_Out, channel64_Kernel61_Valid_Out;

	assign add_kernel61=channel1_Kernel61_Valid_Out & channel2_Kernel61_Valid_Out & channel3_Kernel61_Valid_Out & channel4_Kernel61_Valid_Out & channel5_Kernel61_Valid_Out & channel6_Kernel61_Valid_Out & channel7_Kernel61_Valid_Out & channel8_Kernel61_Valid_Out & channel9_Kernel61_Valid_Out & channel10_Kernel61_Valid_Out & channel11_Kernel61_Valid_Out & channel12_Kernel61_Valid_Out & channel13_Kernel61_Valid_Out & channel14_Kernel61_Valid_Out & channel15_Kernel61_Valid_Out & channel16_Kernel61_Valid_Out & channel17_Kernel61_Valid_Out & channel18_Kernel61_Valid_Out & channel19_Kernel61_Valid_Out & channel20_Kernel61_Valid_Out & channel21_Kernel61_Valid_Out & channel22_Kernel61_Valid_Out & channel23_Kernel61_Valid_Out & channel24_Kernel61_Valid_Out & channel25_Kernel61_Valid_Out & channel26_Kernel61_Valid_Out & channel27_Kernel61_Valid_Out & channel28_Kernel61_Valid_Out & channel29_Kernel61_Valid_Out & channel30_Kernel61_Valid_Out & channel31_Kernel61_Valid_Out & channel32_Kernel61_Valid_Out & channel33_Kernel61_Valid_Out & channel34_Kernel61_Valid_Out & channel35_Kernel61_Valid_Out & channel36_Kernel61_Valid_Out & channel37_Kernel61_Valid_Out & channel38_Kernel61_Valid_Out & channel39_Kernel61_Valid_Out & channel40_Kernel61_Valid_Out & channel41_Kernel61_Valid_Out & channel42_Kernel61_Valid_Out & channel43_Kernel61_Valid_Out & channel44_Kernel61_Valid_Out & channel45_Kernel61_Valid_Out & channel46_Kernel61_Valid_Out & channel47_Kernel61_Valid_Out & channel48_Kernel61_Valid_Out & channel49_Kernel61_Valid_Out & channel50_Kernel61_Valid_Out & channel51_Kernel61_Valid_Out & channel52_Kernel61_Valid_Out & channel53_Kernel61_Valid_Out & channel54_Kernel61_Valid_Out & channel55_Kernel61_Valid_Out & channel56_Kernel61_Valid_Out & channel57_Kernel61_Valid_Out & channel58_Kernel61_Valid_Out & channel59_Kernel61_Valid_Out & channel60_Kernel61_Valid_Out & channel61_Kernel61_Valid_Out & channel62_Kernel61_Valid_Out & channel63_Kernel61_Valid_Out & channel64_Kernel61_Valid_Out;

	wire channel1_Kernel62_Valid_Out, channel2_Kernel62_Valid_Out, channel3_Kernel62_Valid_Out, channel4_Kernel62_Valid_Out, channel5_Kernel62_Valid_Out, channel6_Kernel62_Valid_Out, channel7_Kernel62_Valid_Out, channel8_Kernel62_Valid_Out, channel9_Kernel62_Valid_Out, channel10_Kernel62_Valid_Out, channel11_Kernel62_Valid_Out, channel12_Kernel62_Valid_Out, channel13_Kernel62_Valid_Out, channel14_Kernel62_Valid_Out, channel15_Kernel62_Valid_Out, channel16_Kernel62_Valid_Out, channel17_Kernel62_Valid_Out, channel18_Kernel62_Valid_Out, channel19_Kernel62_Valid_Out, channel20_Kernel62_Valid_Out, channel21_Kernel62_Valid_Out, channel22_Kernel62_Valid_Out, channel23_Kernel62_Valid_Out, channel24_Kernel62_Valid_Out, channel25_Kernel62_Valid_Out, channel26_Kernel62_Valid_Out, channel27_Kernel62_Valid_Out, channel28_Kernel62_Valid_Out, channel29_Kernel62_Valid_Out, channel30_Kernel62_Valid_Out, channel31_Kernel62_Valid_Out, channel32_Kernel62_Valid_Out, channel33_Kernel62_Valid_Out, channel34_Kernel62_Valid_Out, channel35_Kernel62_Valid_Out, channel36_Kernel62_Valid_Out, channel37_Kernel62_Valid_Out, channel38_Kernel62_Valid_Out, channel39_Kernel62_Valid_Out, channel40_Kernel62_Valid_Out, channel41_Kernel62_Valid_Out, channel42_Kernel62_Valid_Out, channel43_Kernel62_Valid_Out, channel44_Kernel62_Valid_Out, channel45_Kernel62_Valid_Out, channel46_Kernel62_Valid_Out, channel47_Kernel62_Valid_Out, channel48_Kernel62_Valid_Out, channel49_Kernel62_Valid_Out, channel50_Kernel62_Valid_Out, channel51_Kernel62_Valid_Out, channel52_Kernel62_Valid_Out, channel53_Kernel62_Valid_Out, channel54_Kernel62_Valid_Out, channel55_Kernel62_Valid_Out, channel56_Kernel62_Valid_Out, channel57_Kernel62_Valid_Out, channel58_Kernel62_Valid_Out, channel59_Kernel62_Valid_Out, channel60_Kernel62_Valid_Out, channel61_Kernel62_Valid_Out, channel62_Kernel62_Valid_Out, channel63_Kernel62_Valid_Out, channel64_Kernel62_Valid_Out;

	assign add_kernel62=channel1_Kernel62_Valid_Out & channel2_Kernel62_Valid_Out & channel3_Kernel62_Valid_Out & channel4_Kernel62_Valid_Out & channel5_Kernel62_Valid_Out & channel6_Kernel62_Valid_Out & channel7_Kernel62_Valid_Out & channel8_Kernel62_Valid_Out & channel9_Kernel62_Valid_Out & channel10_Kernel62_Valid_Out & channel11_Kernel62_Valid_Out & channel12_Kernel62_Valid_Out & channel13_Kernel62_Valid_Out & channel14_Kernel62_Valid_Out & channel15_Kernel62_Valid_Out & channel16_Kernel62_Valid_Out & channel17_Kernel62_Valid_Out & channel18_Kernel62_Valid_Out & channel19_Kernel62_Valid_Out & channel20_Kernel62_Valid_Out & channel21_Kernel62_Valid_Out & channel22_Kernel62_Valid_Out & channel23_Kernel62_Valid_Out & channel24_Kernel62_Valid_Out & channel25_Kernel62_Valid_Out & channel26_Kernel62_Valid_Out & channel27_Kernel62_Valid_Out & channel28_Kernel62_Valid_Out & channel29_Kernel62_Valid_Out & channel30_Kernel62_Valid_Out & channel31_Kernel62_Valid_Out & channel32_Kernel62_Valid_Out & channel33_Kernel62_Valid_Out & channel34_Kernel62_Valid_Out & channel35_Kernel62_Valid_Out & channel36_Kernel62_Valid_Out & channel37_Kernel62_Valid_Out & channel38_Kernel62_Valid_Out & channel39_Kernel62_Valid_Out & channel40_Kernel62_Valid_Out & channel41_Kernel62_Valid_Out & channel42_Kernel62_Valid_Out & channel43_Kernel62_Valid_Out & channel44_Kernel62_Valid_Out & channel45_Kernel62_Valid_Out & channel46_Kernel62_Valid_Out & channel47_Kernel62_Valid_Out & channel48_Kernel62_Valid_Out & channel49_Kernel62_Valid_Out & channel50_Kernel62_Valid_Out & channel51_Kernel62_Valid_Out & channel52_Kernel62_Valid_Out & channel53_Kernel62_Valid_Out & channel54_Kernel62_Valid_Out & channel55_Kernel62_Valid_Out & channel56_Kernel62_Valid_Out & channel57_Kernel62_Valid_Out & channel58_Kernel62_Valid_Out & channel59_Kernel62_Valid_Out & channel60_Kernel62_Valid_Out & channel61_Kernel62_Valid_Out & channel62_Kernel62_Valid_Out & channel63_Kernel62_Valid_Out & channel64_Kernel62_Valid_Out;

	wire channel1_Kernel63_Valid_Out, channel2_Kernel63_Valid_Out, channel3_Kernel63_Valid_Out, channel4_Kernel63_Valid_Out, channel5_Kernel63_Valid_Out, channel6_Kernel63_Valid_Out, channel7_Kernel63_Valid_Out, channel8_Kernel63_Valid_Out, channel9_Kernel63_Valid_Out, channel10_Kernel63_Valid_Out, channel11_Kernel63_Valid_Out, channel12_Kernel63_Valid_Out, channel13_Kernel63_Valid_Out, channel14_Kernel63_Valid_Out, channel15_Kernel63_Valid_Out, channel16_Kernel63_Valid_Out, channel17_Kernel63_Valid_Out, channel18_Kernel63_Valid_Out, channel19_Kernel63_Valid_Out, channel20_Kernel63_Valid_Out, channel21_Kernel63_Valid_Out, channel22_Kernel63_Valid_Out, channel23_Kernel63_Valid_Out, channel24_Kernel63_Valid_Out, channel25_Kernel63_Valid_Out, channel26_Kernel63_Valid_Out, channel27_Kernel63_Valid_Out, channel28_Kernel63_Valid_Out, channel29_Kernel63_Valid_Out, channel30_Kernel63_Valid_Out, channel31_Kernel63_Valid_Out, channel32_Kernel63_Valid_Out, channel33_Kernel63_Valid_Out, channel34_Kernel63_Valid_Out, channel35_Kernel63_Valid_Out, channel36_Kernel63_Valid_Out, channel37_Kernel63_Valid_Out, channel38_Kernel63_Valid_Out, channel39_Kernel63_Valid_Out, channel40_Kernel63_Valid_Out, channel41_Kernel63_Valid_Out, channel42_Kernel63_Valid_Out, channel43_Kernel63_Valid_Out, channel44_Kernel63_Valid_Out, channel45_Kernel63_Valid_Out, channel46_Kernel63_Valid_Out, channel47_Kernel63_Valid_Out, channel48_Kernel63_Valid_Out, channel49_Kernel63_Valid_Out, channel50_Kernel63_Valid_Out, channel51_Kernel63_Valid_Out, channel52_Kernel63_Valid_Out, channel53_Kernel63_Valid_Out, channel54_Kernel63_Valid_Out, channel55_Kernel63_Valid_Out, channel56_Kernel63_Valid_Out, channel57_Kernel63_Valid_Out, channel58_Kernel63_Valid_Out, channel59_Kernel63_Valid_Out, channel60_Kernel63_Valid_Out, channel61_Kernel63_Valid_Out, channel62_Kernel63_Valid_Out, channel63_Kernel63_Valid_Out, channel64_Kernel63_Valid_Out;

	assign add_kernel63=channel1_Kernel63_Valid_Out & channel2_Kernel63_Valid_Out & channel3_Kernel63_Valid_Out & channel4_Kernel63_Valid_Out & channel5_Kernel63_Valid_Out & channel6_Kernel63_Valid_Out & channel7_Kernel63_Valid_Out & channel8_Kernel63_Valid_Out & channel9_Kernel63_Valid_Out & channel10_Kernel63_Valid_Out & channel11_Kernel63_Valid_Out & channel12_Kernel63_Valid_Out & channel13_Kernel63_Valid_Out & channel14_Kernel63_Valid_Out & channel15_Kernel63_Valid_Out & channel16_Kernel63_Valid_Out & channel17_Kernel63_Valid_Out & channel18_Kernel63_Valid_Out & channel19_Kernel63_Valid_Out & channel20_Kernel63_Valid_Out & channel21_Kernel63_Valid_Out & channel22_Kernel63_Valid_Out & channel23_Kernel63_Valid_Out & channel24_Kernel63_Valid_Out & channel25_Kernel63_Valid_Out & channel26_Kernel63_Valid_Out & channel27_Kernel63_Valid_Out & channel28_Kernel63_Valid_Out & channel29_Kernel63_Valid_Out & channel30_Kernel63_Valid_Out & channel31_Kernel63_Valid_Out & channel32_Kernel63_Valid_Out & channel33_Kernel63_Valid_Out & channel34_Kernel63_Valid_Out & channel35_Kernel63_Valid_Out & channel36_Kernel63_Valid_Out & channel37_Kernel63_Valid_Out & channel38_Kernel63_Valid_Out & channel39_Kernel63_Valid_Out & channel40_Kernel63_Valid_Out & channel41_Kernel63_Valid_Out & channel42_Kernel63_Valid_Out & channel43_Kernel63_Valid_Out & channel44_Kernel63_Valid_Out & channel45_Kernel63_Valid_Out & channel46_Kernel63_Valid_Out & channel47_Kernel63_Valid_Out & channel48_Kernel63_Valid_Out & channel49_Kernel63_Valid_Out & channel50_Kernel63_Valid_Out & channel51_Kernel63_Valid_Out & channel52_Kernel63_Valid_Out & channel53_Kernel63_Valid_Out & channel54_Kernel63_Valid_Out & channel55_Kernel63_Valid_Out & channel56_Kernel63_Valid_Out & channel57_Kernel63_Valid_Out & channel58_Kernel63_Valid_Out & channel59_Kernel63_Valid_Out & channel60_Kernel63_Valid_Out & channel61_Kernel63_Valid_Out & channel62_Kernel63_Valid_Out & channel63_Kernel63_Valid_Out & channel64_Kernel63_Valid_Out;

	wire channel1_Kernel64_Valid_Out, channel2_Kernel64_Valid_Out, channel3_Kernel64_Valid_Out, channel4_Kernel64_Valid_Out, channel5_Kernel64_Valid_Out, channel6_Kernel64_Valid_Out, channel7_Kernel64_Valid_Out, channel8_Kernel64_Valid_Out, channel9_Kernel64_Valid_Out, channel10_Kernel64_Valid_Out, channel11_Kernel64_Valid_Out, channel12_Kernel64_Valid_Out, channel13_Kernel64_Valid_Out, channel14_Kernel64_Valid_Out, channel15_Kernel64_Valid_Out, channel16_Kernel64_Valid_Out, channel17_Kernel64_Valid_Out, channel18_Kernel64_Valid_Out, channel19_Kernel64_Valid_Out, channel20_Kernel64_Valid_Out, channel21_Kernel64_Valid_Out, channel22_Kernel64_Valid_Out, channel23_Kernel64_Valid_Out, channel24_Kernel64_Valid_Out, channel25_Kernel64_Valid_Out, channel26_Kernel64_Valid_Out, channel27_Kernel64_Valid_Out, channel28_Kernel64_Valid_Out, channel29_Kernel64_Valid_Out, channel30_Kernel64_Valid_Out, channel31_Kernel64_Valid_Out, channel32_Kernel64_Valid_Out, channel33_Kernel64_Valid_Out, channel34_Kernel64_Valid_Out, channel35_Kernel64_Valid_Out, channel36_Kernel64_Valid_Out, channel37_Kernel64_Valid_Out, channel38_Kernel64_Valid_Out, channel39_Kernel64_Valid_Out, channel40_Kernel64_Valid_Out, channel41_Kernel64_Valid_Out, channel42_Kernel64_Valid_Out, channel43_Kernel64_Valid_Out, channel44_Kernel64_Valid_Out, channel45_Kernel64_Valid_Out, channel46_Kernel64_Valid_Out, channel47_Kernel64_Valid_Out, channel48_Kernel64_Valid_Out, channel49_Kernel64_Valid_Out, channel50_Kernel64_Valid_Out, channel51_Kernel64_Valid_Out, channel52_Kernel64_Valid_Out, channel53_Kernel64_Valid_Out, channel54_Kernel64_Valid_Out, channel55_Kernel64_Valid_Out, channel56_Kernel64_Valid_Out, channel57_Kernel64_Valid_Out, channel58_Kernel64_Valid_Out, channel59_Kernel64_Valid_Out, channel60_Kernel64_Valid_Out, channel61_Kernel64_Valid_Out, channel62_Kernel64_Valid_Out, channel63_Kernel64_Valid_Out, channel64_Kernel64_Valid_Out;

	assign add_kernel64=channel1_Kernel64_Valid_Out & channel2_Kernel64_Valid_Out & channel3_Kernel64_Valid_Out & channel4_Kernel64_Valid_Out & channel5_Kernel64_Valid_Out & channel6_Kernel64_Valid_Out & channel7_Kernel64_Valid_Out & channel8_Kernel64_Valid_Out & channel9_Kernel64_Valid_Out & channel10_Kernel64_Valid_Out & channel11_Kernel64_Valid_Out & channel12_Kernel64_Valid_Out & channel13_Kernel64_Valid_Out & channel14_Kernel64_Valid_Out & channel15_Kernel64_Valid_Out & channel16_Kernel64_Valid_Out & channel17_Kernel64_Valid_Out & channel18_Kernel64_Valid_Out & channel19_Kernel64_Valid_Out & channel20_Kernel64_Valid_Out & channel21_Kernel64_Valid_Out & channel22_Kernel64_Valid_Out & channel23_Kernel64_Valid_Out & channel24_Kernel64_Valid_Out & channel25_Kernel64_Valid_Out & channel26_Kernel64_Valid_Out & channel27_Kernel64_Valid_Out & channel28_Kernel64_Valid_Out & channel29_Kernel64_Valid_Out & channel30_Kernel64_Valid_Out & channel31_Kernel64_Valid_Out & channel32_Kernel64_Valid_Out & channel33_Kernel64_Valid_Out & channel34_Kernel64_Valid_Out & channel35_Kernel64_Valid_Out & channel36_Kernel64_Valid_Out & channel37_Kernel64_Valid_Out & channel38_Kernel64_Valid_Out & channel39_Kernel64_Valid_Out & channel40_Kernel64_Valid_Out & channel41_Kernel64_Valid_Out & channel42_Kernel64_Valid_Out & channel43_Kernel64_Valid_Out & channel44_Kernel64_Valid_Out & channel45_Kernel64_Valid_Out & channel46_Kernel64_Valid_Out & channel47_Kernel64_Valid_Out & channel48_Kernel64_Valid_Out & channel49_Kernel64_Valid_Out & channel50_Kernel64_Valid_Out & channel51_Kernel64_Valid_Out & channel52_Kernel64_Valid_Out & channel53_Kernel64_Valid_Out & channel54_Kernel64_Valid_Out & channel55_Kernel64_Valid_Out & channel56_Kernel64_Valid_Out & channel57_Kernel64_Valid_Out & channel58_Kernel64_Valid_Out & channel59_Kernel64_Valid_Out & channel60_Kernel64_Valid_Out & channel61_Kernel64_Valid_Out & channel62_Kernel64_Valid_Out & channel63_Kernel64_Valid_Out & channel64_Kernel64_Valid_Out;

	wire channel1_Kernel65_Valid_Out, channel2_Kernel65_Valid_Out, channel3_Kernel65_Valid_Out, channel4_Kernel65_Valid_Out, channel5_Kernel65_Valid_Out, channel6_Kernel65_Valid_Out, channel7_Kernel65_Valid_Out, channel8_Kernel65_Valid_Out, channel9_Kernel65_Valid_Out, channel10_Kernel65_Valid_Out, channel11_Kernel65_Valid_Out, channel12_Kernel65_Valid_Out, channel13_Kernel65_Valid_Out, channel14_Kernel65_Valid_Out, channel15_Kernel65_Valid_Out, channel16_Kernel65_Valid_Out, channel17_Kernel65_Valid_Out, channel18_Kernel65_Valid_Out, channel19_Kernel65_Valid_Out, channel20_Kernel65_Valid_Out, channel21_Kernel65_Valid_Out, channel22_Kernel65_Valid_Out, channel23_Kernel65_Valid_Out, channel24_Kernel65_Valid_Out, channel25_Kernel65_Valid_Out, channel26_Kernel65_Valid_Out, channel27_Kernel65_Valid_Out, channel28_Kernel65_Valid_Out, channel29_Kernel65_Valid_Out, channel30_Kernel65_Valid_Out, channel31_Kernel65_Valid_Out, channel32_Kernel65_Valid_Out, channel33_Kernel65_Valid_Out, channel34_Kernel65_Valid_Out, channel35_Kernel65_Valid_Out, channel36_Kernel65_Valid_Out, channel37_Kernel65_Valid_Out, channel38_Kernel65_Valid_Out, channel39_Kernel65_Valid_Out, channel40_Kernel65_Valid_Out, channel41_Kernel65_Valid_Out, channel42_Kernel65_Valid_Out, channel43_Kernel65_Valid_Out, channel44_Kernel65_Valid_Out, channel45_Kernel65_Valid_Out, channel46_Kernel65_Valid_Out, channel47_Kernel65_Valid_Out, channel48_Kernel65_Valid_Out, channel49_Kernel65_Valid_Out, channel50_Kernel65_Valid_Out, channel51_Kernel65_Valid_Out, channel52_Kernel65_Valid_Out, channel53_Kernel65_Valid_Out, channel54_Kernel65_Valid_Out, channel55_Kernel65_Valid_Out, channel56_Kernel65_Valid_Out, channel57_Kernel65_Valid_Out, channel58_Kernel65_Valid_Out, channel59_Kernel65_Valid_Out, channel60_Kernel65_Valid_Out, channel61_Kernel65_Valid_Out, channel62_Kernel65_Valid_Out, channel63_Kernel65_Valid_Out, channel64_Kernel65_Valid_Out;

	assign add_kernel65=channel1_Kernel65_Valid_Out & channel2_Kernel65_Valid_Out & channel3_Kernel65_Valid_Out & channel4_Kernel65_Valid_Out & channel5_Kernel65_Valid_Out & channel6_Kernel65_Valid_Out & channel7_Kernel65_Valid_Out & channel8_Kernel65_Valid_Out & channel9_Kernel65_Valid_Out & channel10_Kernel65_Valid_Out & channel11_Kernel65_Valid_Out & channel12_Kernel65_Valid_Out & channel13_Kernel65_Valid_Out & channel14_Kernel65_Valid_Out & channel15_Kernel65_Valid_Out & channel16_Kernel65_Valid_Out & channel17_Kernel65_Valid_Out & channel18_Kernel65_Valid_Out & channel19_Kernel65_Valid_Out & channel20_Kernel65_Valid_Out & channel21_Kernel65_Valid_Out & channel22_Kernel65_Valid_Out & channel23_Kernel65_Valid_Out & channel24_Kernel65_Valid_Out & channel25_Kernel65_Valid_Out & channel26_Kernel65_Valid_Out & channel27_Kernel65_Valid_Out & channel28_Kernel65_Valid_Out & channel29_Kernel65_Valid_Out & channel30_Kernel65_Valid_Out & channel31_Kernel65_Valid_Out & channel32_Kernel65_Valid_Out & channel33_Kernel65_Valid_Out & channel34_Kernel65_Valid_Out & channel35_Kernel65_Valid_Out & channel36_Kernel65_Valid_Out & channel37_Kernel65_Valid_Out & channel38_Kernel65_Valid_Out & channel39_Kernel65_Valid_Out & channel40_Kernel65_Valid_Out & channel41_Kernel65_Valid_Out & channel42_Kernel65_Valid_Out & channel43_Kernel65_Valid_Out & channel44_Kernel65_Valid_Out & channel45_Kernel65_Valid_Out & channel46_Kernel65_Valid_Out & channel47_Kernel65_Valid_Out & channel48_Kernel65_Valid_Out & channel49_Kernel65_Valid_Out & channel50_Kernel65_Valid_Out & channel51_Kernel65_Valid_Out & channel52_Kernel65_Valid_Out & channel53_Kernel65_Valid_Out & channel54_Kernel65_Valid_Out & channel55_Kernel65_Valid_Out & channel56_Kernel65_Valid_Out & channel57_Kernel65_Valid_Out & channel58_Kernel65_Valid_Out & channel59_Kernel65_Valid_Out & channel60_Kernel65_Valid_Out & channel61_Kernel65_Valid_Out & channel62_Kernel65_Valid_Out & channel63_Kernel65_Valid_Out & channel64_Kernel65_Valid_Out;

	wire channel1_Kernel66_Valid_Out, channel2_Kernel66_Valid_Out, channel3_Kernel66_Valid_Out, channel4_Kernel66_Valid_Out, channel5_Kernel66_Valid_Out, channel6_Kernel66_Valid_Out, channel7_Kernel66_Valid_Out, channel8_Kernel66_Valid_Out, channel9_Kernel66_Valid_Out, channel10_Kernel66_Valid_Out, channel11_Kernel66_Valid_Out, channel12_Kernel66_Valid_Out, channel13_Kernel66_Valid_Out, channel14_Kernel66_Valid_Out, channel15_Kernel66_Valid_Out, channel16_Kernel66_Valid_Out, channel17_Kernel66_Valid_Out, channel18_Kernel66_Valid_Out, channel19_Kernel66_Valid_Out, channel20_Kernel66_Valid_Out, channel21_Kernel66_Valid_Out, channel22_Kernel66_Valid_Out, channel23_Kernel66_Valid_Out, channel24_Kernel66_Valid_Out, channel25_Kernel66_Valid_Out, channel26_Kernel66_Valid_Out, channel27_Kernel66_Valid_Out, channel28_Kernel66_Valid_Out, channel29_Kernel66_Valid_Out, channel30_Kernel66_Valid_Out, channel31_Kernel66_Valid_Out, channel32_Kernel66_Valid_Out, channel33_Kernel66_Valid_Out, channel34_Kernel66_Valid_Out, channel35_Kernel66_Valid_Out, channel36_Kernel66_Valid_Out, channel37_Kernel66_Valid_Out, channel38_Kernel66_Valid_Out, channel39_Kernel66_Valid_Out, channel40_Kernel66_Valid_Out, channel41_Kernel66_Valid_Out, channel42_Kernel66_Valid_Out, channel43_Kernel66_Valid_Out, channel44_Kernel66_Valid_Out, channel45_Kernel66_Valid_Out, channel46_Kernel66_Valid_Out, channel47_Kernel66_Valid_Out, channel48_Kernel66_Valid_Out, channel49_Kernel66_Valid_Out, channel50_Kernel66_Valid_Out, channel51_Kernel66_Valid_Out, channel52_Kernel66_Valid_Out, channel53_Kernel66_Valid_Out, channel54_Kernel66_Valid_Out, channel55_Kernel66_Valid_Out, channel56_Kernel66_Valid_Out, channel57_Kernel66_Valid_Out, channel58_Kernel66_Valid_Out, channel59_Kernel66_Valid_Out, channel60_Kernel66_Valid_Out, channel61_Kernel66_Valid_Out, channel62_Kernel66_Valid_Out, channel63_Kernel66_Valid_Out, channel64_Kernel66_Valid_Out;

	assign add_kernel66=channel1_Kernel66_Valid_Out & channel2_Kernel66_Valid_Out & channel3_Kernel66_Valid_Out & channel4_Kernel66_Valid_Out & channel5_Kernel66_Valid_Out & channel6_Kernel66_Valid_Out & channel7_Kernel66_Valid_Out & channel8_Kernel66_Valid_Out & channel9_Kernel66_Valid_Out & channel10_Kernel66_Valid_Out & channel11_Kernel66_Valid_Out & channel12_Kernel66_Valid_Out & channel13_Kernel66_Valid_Out & channel14_Kernel66_Valid_Out & channel15_Kernel66_Valid_Out & channel16_Kernel66_Valid_Out & channel17_Kernel66_Valid_Out & channel18_Kernel66_Valid_Out & channel19_Kernel66_Valid_Out & channel20_Kernel66_Valid_Out & channel21_Kernel66_Valid_Out & channel22_Kernel66_Valid_Out & channel23_Kernel66_Valid_Out & channel24_Kernel66_Valid_Out & channel25_Kernel66_Valid_Out & channel26_Kernel66_Valid_Out & channel27_Kernel66_Valid_Out & channel28_Kernel66_Valid_Out & channel29_Kernel66_Valid_Out & channel30_Kernel66_Valid_Out & channel31_Kernel66_Valid_Out & channel32_Kernel66_Valid_Out & channel33_Kernel66_Valid_Out & channel34_Kernel66_Valid_Out & channel35_Kernel66_Valid_Out & channel36_Kernel66_Valid_Out & channel37_Kernel66_Valid_Out & channel38_Kernel66_Valid_Out & channel39_Kernel66_Valid_Out & channel40_Kernel66_Valid_Out & channel41_Kernel66_Valid_Out & channel42_Kernel66_Valid_Out & channel43_Kernel66_Valid_Out & channel44_Kernel66_Valid_Out & channel45_Kernel66_Valid_Out & channel46_Kernel66_Valid_Out & channel47_Kernel66_Valid_Out & channel48_Kernel66_Valid_Out & channel49_Kernel66_Valid_Out & channel50_Kernel66_Valid_Out & channel51_Kernel66_Valid_Out & channel52_Kernel66_Valid_Out & channel53_Kernel66_Valid_Out & channel54_Kernel66_Valid_Out & channel55_Kernel66_Valid_Out & channel56_Kernel66_Valid_Out & channel57_Kernel66_Valid_Out & channel58_Kernel66_Valid_Out & channel59_Kernel66_Valid_Out & channel60_Kernel66_Valid_Out & channel61_Kernel66_Valid_Out & channel62_Kernel66_Valid_Out & channel63_Kernel66_Valid_Out & channel64_Kernel66_Valid_Out;

	wire channel1_Kernel67_Valid_Out, channel2_Kernel67_Valid_Out, channel3_Kernel67_Valid_Out, channel4_Kernel67_Valid_Out, channel5_Kernel67_Valid_Out, channel6_Kernel67_Valid_Out, channel7_Kernel67_Valid_Out, channel8_Kernel67_Valid_Out, channel9_Kernel67_Valid_Out, channel10_Kernel67_Valid_Out, channel11_Kernel67_Valid_Out, channel12_Kernel67_Valid_Out, channel13_Kernel67_Valid_Out, channel14_Kernel67_Valid_Out, channel15_Kernel67_Valid_Out, channel16_Kernel67_Valid_Out, channel17_Kernel67_Valid_Out, channel18_Kernel67_Valid_Out, channel19_Kernel67_Valid_Out, channel20_Kernel67_Valid_Out, channel21_Kernel67_Valid_Out, channel22_Kernel67_Valid_Out, channel23_Kernel67_Valid_Out, channel24_Kernel67_Valid_Out, channel25_Kernel67_Valid_Out, channel26_Kernel67_Valid_Out, channel27_Kernel67_Valid_Out, channel28_Kernel67_Valid_Out, channel29_Kernel67_Valid_Out, channel30_Kernel67_Valid_Out, channel31_Kernel67_Valid_Out, channel32_Kernel67_Valid_Out, channel33_Kernel67_Valid_Out, channel34_Kernel67_Valid_Out, channel35_Kernel67_Valid_Out, channel36_Kernel67_Valid_Out, channel37_Kernel67_Valid_Out, channel38_Kernel67_Valid_Out, channel39_Kernel67_Valid_Out, channel40_Kernel67_Valid_Out, channel41_Kernel67_Valid_Out, channel42_Kernel67_Valid_Out, channel43_Kernel67_Valid_Out, channel44_Kernel67_Valid_Out, channel45_Kernel67_Valid_Out, channel46_Kernel67_Valid_Out, channel47_Kernel67_Valid_Out, channel48_Kernel67_Valid_Out, channel49_Kernel67_Valid_Out, channel50_Kernel67_Valid_Out, channel51_Kernel67_Valid_Out, channel52_Kernel67_Valid_Out, channel53_Kernel67_Valid_Out, channel54_Kernel67_Valid_Out, channel55_Kernel67_Valid_Out, channel56_Kernel67_Valid_Out, channel57_Kernel67_Valid_Out, channel58_Kernel67_Valid_Out, channel59_Kernel67_Valid_Out, channel60_Kernel67_Valid_Out, channel61_Kernel67_Valid_Out, channel62_Kernel67_Valid_Out, channel63_Kernel67_Valid_Out, channel64_Kernel67_Valid_Out;

	assign add_kernel67=channel1_Kernel67_Valid_Out & channel2_Kernel67_Valid_Out & channel3_Kernel67_Valid_Out & channel4_Kernel67_Valid_Out & channel5_Kernel67_Valid_Out & channel6_Kernel67_Valid_Out & channel7_Kernel67_Valid_Out & channel8_Kernel67_Valid_Out & channel9_Kernel67_Valid_Out & channel10_Kernel67_Valid_Out & channel11_Kernel67_Valid_Out & channel12_Kernel67_Valid_Out & channel13_Kernel67_Valid_Out & channel14_Kernel67_Valid_Out & channel15_Kernel67_Valid_Out & channel16_Kernel67_Valid_Out & channel17_Kernel67_Valid_Out & channel18_Kernel67_Valid_Out & channel19_Kernel67_Valid_Out & channel20_Kernel67_Valid_Out & channel21_Kernel67_Valid_Out & channel22_Kernel67_Valid_Out & channel23_Kernel67_Valid_Out & channel24_Kernel67_Valid_Out & channel25_Kernel67_Valid_Out & channel26_Kernel67_Valid_Out & channel27_Kernel67_Valid_Out & channel28_Kernel67_Valid_Out & channel29_Kernel67_Valid_Out & channel30_Kernel67_Valid_Out & channel31_Kernel67_Valid_Out & channel32_Kernel67_Valid_Out & channel33_Kernel67_Valid_Out & channel34_Kernel67_Valid_Out & channel35_Kernel67_Valid_Out & channel36_Kernel67_Valid_Out & channel37_Kernel67_Valid_Out & channel38_Kernel67_Valid_Out & channel39_Kernel67_Valid_Out & channel40_Kernel67_Valid_Out & channel41_Kernel67_Valid_Out & channel42_Kernel67_Valid_Out & channel43_Kernel67_Valid_Out & channel44_Kernel67_Valid_Out & channel45_Kernel67_Valid_Out & channel46_Kernel67_Valid_Out & channel47_Kernel67_Valid_Out & channel48_Kernel67_Valid_Out & channel49_Kernel67_Valid_Out & channel50_Kernel67_Valid_Out & channel51_Kernel67_Valid_Out & channel52_Kernel67_Valid_Out & channel53_Kernel67_Valid_Out & channel54_Kernel67_Valid_Out & channel55_Kernel67_Valid_Out & channel56_Kernel67_Valid_Out & channel57_Kernel67_Valid_Out & channel58_Kernel67_Valid_Out & channel59_Kernel67_Valid_Out & channel60_Kernel67_Valid_Out & channel61_Kernel67_Valid_Out & channel62_Kernel67_Valid_Out & channel63_Kernel67_Valid_Out & channel64_Kernel67_Valid_Out;

	wire channel1_Kernel68_Valid_Out, channel2_Kernel68_Valid_Out, channel3_Kernel68_Valid_Out, channel4_Kernel68_Valid_Out, channel5_Kernel68_Valid_Out, channel6_Kernel68_Valid_Out, channel7_Kernel68_Valid_Out, channel8_Kernel68_Valid_Out, channel9_Kernel68_Valid_Out, channel10_Kernel68_Valid_Out, channel11_Kernel68_Valid_Out, channel12_Kernel68_Valid_Out, channel13_Kernel68_Valid_Out, channel14_Kernel68_Valid_Out, channel15_Kernel68_Valid_Out, channel16_Kernel68_Valid_Out, channel17_Kernel68_Valid_Out, channel18_Kernel68_Valid_Out, channel19_Kernel68_Valid_Out, channel20_Kernel68_Valid_Out, channel21_Kernel68_Valid_Out, channel22_Kernel68_Valid_Out, channel23_Kernel68_Valid_Out, channel24_Kernel68_Valid_Out, channel25_Kernel68_Valid_Out, channel26_Kernel68_Valid_Out, channel27_Kernel68_Valid_Out, channel28_Kernel68_Valid_Out, channel29_Kernel68_Valid_Out, channel30_Kernel68_Valid_Out, channel31_Kernel68_Valid_Out, channel32_Kernel68_Valid_Out, channel33_Kernel68_Valid_Out, channel34_Kernel68_Valid_Out, channel35_Kernel68_Valid_Out, channel36_Kernel68_Valid_Out, channel37_Kernel68_Valid_Out, channel38_Kernel68_Valid_Out, channel39_Kernel68_Valid_Out, channel40_Kernel68_Valid_Out, channel41_Kernel68_Valid_Out, channel42_Kernel68_Valid_Out, channel43_Kernel68_Valid_Out, channel44_Kernel68_Valid_Out, channel45_Kernel68_Valid_Out, channel46_Kernel68_Valid_Out, channel47_Kernel68_Valid_Out, channel48_Kernel68_Valid_Out, channel49_Kernel68_Valid_Out, channel50_Kernel68_Valid_Out, channel51_Kernel68_Valid_Out, channel52_Kernel68_Valid_Out, channel53_Kernel68_Valid_Out, channel54_Kernel68_Valid_Out, channel55_Kernel68_Valid_Out, channel56_Kernel68_Valid_Out, channel57_Kernel68_Valid_Out, channel58_Kernel68_Valid_Out, channel59_Kernel68_Valid_Out, channel60_Kernel68_Valid_Out, channel61_Kernel68_Valid_Out, channel62_Kernel68_Valid_Out, channel63_Kernel68_Valid_Out, channel64_Kernel68_Valid_Out;

	assign add_kernel68=channel1_Kernel68_Valid_Out & channel2_Kernel68_Valid_Out & channel3_Kernel68_Valid_Out & channel4_Kernel68_Valid_Out & channel5_Kernel68_Valid_Out & channel6_Kernel68_Valid_Out & channel7_Kernel68_Valid_Out & channel8_Kernel68_Valid_Out & channel9_Kernel68_Valid_Out & channel10_Kernel68_Valid_Out & channel11_Kernel68_Valid_Out & channel12_Kernel68_Valid_Out & channel13_Kernel68_Valid_Out & channel14_Kernel68_Valid_Out & channel15_Kernel68_Valid_Out & channel16_Kernel68_Valid_Out & channel17_Kernel68_Valid_Out & channel18_Kernel68_Valid_Out & channel19_Kernel68_Valid_Out & channel20_Kernel68_Valid_Out & channel21_Kernel68_Valid_Out & channel22_Kernel68_Valid_Out & channel23_Kernel68_Valid_Out & channel24_Kernel68_Valid_Out & channel25_Kernel68_Valid_Out & channel26_Kernel68_Valid_Out & channel27_Kernel68_Valid_Out & channel28_Kernel68_Valid_Out & channel29_Kernel68_Valid_Out & channel30_Kernel68_Valid_Out & channel31_Kernel68_Valid_Out & channel32_Kernel68_Valid_Out & channel33_Kernel68_Valid_Out & channel34_Kernel68_Valid_Out & channel35_Kernel68_Valid_Out & channel36_Kernel68_Valid_Out & channel37_Kernel68_Valid_Out & channel38_Kernel68_Valid_Out & channel39_Kernel68_Valid_Out & channel40_Kernel68_Valid_Out & channel41_Kernel68_Valid_Out & channel42_Kernel68_Valid_Out & channel43_Kernel68_Valid_Out & channel44_Kernel68_Valid_Out & channel45_Kernel68_Valid_Out & channel46_Kernel68_Valid_Out & channel47_Kernel68_Valid_Out & channel48_Kernel68_Valid_Out & channel49_Kernel68_Valid_Out & channel50_Kernel68_Valid_Out & channel51_Kernel68_Valid_Out & channel52_Kernel68_Valid_Out & channel53_Kernel68_Valid_Out & channel54_Kernel68_Valid_Out & channel55_Kernel68_Valid_Out & channel56_Kernel68_Valid_Out & channel57_Kernel68_Valid_Out & channel58_Kernel68_Valid_Out & channel59_Kernel68_Valid_Out & channel60_Kernel68_Valid_Out & channel61_Kernel68_Valid_Out & channel62_Kernel68_Valid_Out & channel63_Kernel68_Valid_Out & channel64_Kernel68_Valid_Out;

	wire channel1_Kernel69_Valid_Out, channel2_Kernel69_Valid_Out, channel3_Kernel69_Valid_Out, channel4_Kernel69_Valid_Out, channel5_Kernel69_Valid_Out, channel6_Kernel69_Valid_Out, channel7_Kernel69_Valid_Out, channel8_Kernel69_Valid_Out, channel9_Kernel69_Valid_Out, channel10_Kernel69_Valid_Out, channel11_Kernel69_Valid_Out, channel12_Kernel69_Valid_Out, channel13_Kernel69_Valid_Out, channel14_Kernel69_Valid_Out, channel15_Kernel69_Valid_Out, channel16_Kernel69_Valid_Out, channel17_Kernel69_Valid_Out, channel18_Kernel69_Valid_Out, channel19_Kernel69_Valid_Out, channel20_Kernel69_Valid_Out, channel21_Kernel69_Valid_Out, channel22_Kernel69_Valid_Out, channel23_Kernel69_Valid_Out, channel24_Kernel69_Valid_Out, channel25_Kernel69_Valid_Out, channel26_Kernel69_Valid_Out, channel27_Kernel69_Valid_Out, channel28_Kernel69_Valid_Out, channel29_Kernel69_Valid_Out, channel30_Kernel69_Valid_Out, channel31_Kernel69_Valid_Out, channel32_Kernel69_Valid_Out, channel33_Kernel69_Valid_Out, channel34_Kernel69_Valid_Out, channel35_Kernel69_Valid_Out, channel36_Kernel69_Valid_Out, channel37_Kernel69_Valid_Out, channel38_Kernel69_Valid_Out, channel39_Kernel69_Valid_Out, channel40_Kernel69_Valid_Out, channel41_Kernel69_Valid_Out, channel42_Kernel69_Valid_Out, channel43_Kernel69_Valid_Out, channel44_Kernel69_Valid_Out, channel45_Kernel69_Valid_Out, channel46_Kernel69_Valid_Out, channel47_Kernel69_Valid_Out, channel48_Kernel69_Valid_Out, channel49_Kernel69_Valid_Out, channel50_Kernel69_Valid_Out, channel51_Kernel69_Valid_Out, channel52_Kernel69_Valid_Out, channel53_Kernel69_Valid_Out, channel54_Kernel69_Valid_Out, channel55_Kernel69_Valid_Out, channel56_Kernel69_Valid_Out, channel57_Kernel69_Valid_Out, channel58_Kernel69_Valid_Out, channel59_Kernel69_Valid_Out, channel60_Kernel69_Valid_Out, channel61_Kernel69_Valid_Out, channel62_Kernel69_Valid_Out, channel63_Kernel69_Valid_Out, channel64_Kernel69_Valid_Out;

	assign add_kernel69=channel1_Kernel69_Valid_Out & channel2_Kernel69_Valid_Out & channel3_Kernel69_Valid_Out & channel4_Kernel69_Valid_Out & channel5_Kernel69_Valid_Out & channel6_Kernel69_Valid_Out & channel7_Kernel69_Valid_Out & channel8_Kernel69_Valid_Out & channel9_Kernel69_Valid_Out & channel10_Kernel69_Valid_Out & channel11_Kernel69_Valid_Out & channel12_Kernel69_Valid_Out & channel13_Kernel69_Valid_Out & channel14_Kernel69_Valid_Out & channel15_Kernel69_Valid_Out & channel16_Kernel69_Valid_Out & channel17_Kernel69_Valid_Out & channel18_Kernel69_Valid_Out & channel19_Kernel69_Valid_Out & channel20_Kernel69_Valid_Out & channel21_Kernel69_Valid_Out & channel22_Kernel69_Valid_Out & channel23_Kernel69_Valid_Out & channel24_Kernel69_Valid_Out & channel25_Kernel69_Valid_Out & channel26_Kernel69_Valid_Out & channel27_Kernel69_Valid_Out & channel28_Kernel69_Valid_Out & channel29_Kernel69_Valid_Out & channel30_Kernel69_Valid_Out & channel31_Kernel69_Valid_Out & channel32_Kernel69_Valid_Out & channel33_Kernel69_Valid_Out & channel34_Kernel69_Valid_Out & channel35_Kernel69_Valid_Out & channel36_Kernel69_Valid_Out & channel37_Kernel69_Valid_Out & channel38_Kernel69_Valid_Out & channel39_Kernel69_Valid_Out & channel40_Kernel69_Valid_Out & channel41_Kernel69_Valid_Out & channel42_Kernel69_Valid_Out & channel43_Kernel69_Valid_Out & channel44_Kernel69_Valid_Out & channel45_Kernel69_Valid_Out & channel46_Kernel69_Valid_Out & channel47_Kernel69_Valid_Out & channel48_Kernel69_Valid_Out & channel49_Kernel69_Valid_Out & channel50_Kernel69_Valid_Out & channel51_Kernel69_Valid_Out & channel52_Kernel69_Valid_Out & channel53_Kernel69_Valid_Out & channel54_Kernel69_Valid_Out & channel55_Kernel69_Valid_Out & channel56_Kernel69_Valid_Out & channel57_Kernel69_Valid_Out & channel58_Kernel69_Valid_Out & channel59_Kernel69_Valid_Out & channel60_Kernel69_Valid_Out & channel61_Kernel69_Valid_Out & channel62_Kernel69_Valid_Out & channel63_Kernel69_Valid_Out & channel64_Kernel69_Valid_Out;

	wire channel1_Kernel70_Valid_Out, channel2_Kernel70_Valid_Out, channel3_Kernel70_Valid_Out, channel4_Kernel70_Valid_Out, channel5_Kernel70_Valid_Out, channel6_Kernel70_Valid_Out, channel7_Kernel70_Valid_Out, channel8_Kernel70_Valid_Out, channel9_Kernel70_Valid_Out, channel10_Kernel70_Valid_Out, channel11_Kernel70_Valid_Out, channel12_Kernel70_Valid_Out, channel13_Kernel70_Valid_Out, channel14_Kernel70_Valid_Out, channel15_Kernel70_Valid_Out, channel16_Kernel70_Valid_Out, channel17_Kernel70_Valid_Out, channel18_Kernel70_Valid_Out, channel19_Kernel70_Valid_Out, channel20_Kernel70_Valid_Out, channel21_Kernel70_Valid_Out, channel22_Kernel70_Valid_Out, channel23_Kernel70_Valid_Out, channel24_Kernel70_Valid_Out, channel25_Kernel70_Valid_Out, channel26_Kernel70_Valid_Out, channel27_Kernel70_Valid_Out, channel28_Kernel70_Valid_Out, channel29_Kernel70_Valid_Out, channel30_Kernel70_Valid_Out, channel31_Kernel70_Valid_Out, channel32_Kernel70_Valid_Out, channel33_Kernel70_Valid_Out, channel34_Kernel70_Valid_Out, channel35_Kernel70_Valid_Out, channel36_Kernel70_Valid_Out, channel37_Kernel70_Valid_Out, channel38_Kernel70_Valid_Out, channel39_Kernel70_Valid_Out, channel40_Kernel70_Valid_Out, channel41_Kernel70_Valid_Out, channel42_Kernel70_Valid_Out, channel43_Kernel70_Valid_Out, channel44_Kernel70_Valid_Out, channel45_Kernel70_Valid_Out, channel46_Kernel70_Valid_Out, channel47_Kernel70_Valid_Out, channel48_Kernel70_Valid_Out, channel49_Kernel70_Valid_Out, channel50_Kernel70_Valid_Out, channel51_Kernel70_Valid_Out, channel52_Kernel70_Valid_Out, channel53_Kernel70_Valid_Out, channel54_Kernel70_Valid_Out, channel55_Kernel70_Valid_Out, channel56_Kernel70_Valid_Out, channel57_Kernel70_Valid_Out, channel58_Kernel70_Valid_Out, channel59_Kernel70_Valid_Out, channel60_Kernel70_Valid_Out, channel61_Kernel70_Valid_Out, channel62_Kernel70_Valid_Out, channel63_Kernel70_Valid_Out, channel64_Kernel70_Valid_Out;

	assign add_kernel70=channel1_Kernel70_Valid_Out & channel2_Kernel70_Valid_Out & channel3_Kernel70_Valid_Out & channel4_Kernel70_Valid_Out & channel5_Kernel70_Valid_Out & channel6_Kernel70_Valid_Out & channel7_Kernel70_Valid_Out & channel8_Kernel70_Valid_Out & channel9_Kernel70_Valid_Out & channel10_Kernel70_Valid_Out & channel11_Kernel70_Valid_Out & channel12_Kernel70_Valid_Out & channel13_Kernel70_Valid_Out & channel14_Kernel70_Valid_Out & channel15_Kernel70_Valid_Out & channel16_Kernel70_Valid_Out & channel17_Kernel70_Valid_Out & channel18_Kernel70_Valid_Out & channel19_Kernel70_Valid_Out & channel20_Kernel70_Valid_Out & channel21_Kernel70_Valid_Out & channel22_Kernel70_Valid_Out & channel23_Kernel70_Valid_Out & channel24_Kernel70_Valid_Out & channel25_Kernel70_Valid_Out & channel26_Kernel70_Valid_Out & channel27_Kernel70_Valid_Out & channel28_Kernel70_Valid_Out & channel29_Kernel70_Valid_Out & channel30_Kernel70_Valid_Out & channel31_Kernel70_Valid_Out & channel32_Kernel70_Valid_Out & channel33_Kernel70_Valid_Out & channel34_Kernel70_Valid_Out & channel35_Kernel70_Valid_Out & channel36_Kernel70_Valid_Out & channel37_Kernel70_Valid_Out & channel38_Kernel70_Valid_Out & channel39_Kernel70_Valid_Out & channel40_Kernel70_Valid_Out & channel41_Kernel70_Valid_Out & channel42_Kernel70_Valid_Out & channel43_Kernel70_Valid_Out & channel44_Kernel70_Valid_Out & channel45_Kernel70_Valid_Out & channel46_Kernel70_Valid_Out & channel47_Kernel70_Valid_Out & channel48_Kernel70_Valid_Out & channel49_Kernel70_Valid_Out & channel50_Kernel70_Valid_Out & channel51_Kernel70_Valid_Out & channel52_Kernel70_Valid_Out & channel53_Kernel70_Valid_Out & channel54_Kernel70_Valid_Out & channel55_Kernel70_Valid_Out & channel56_Kernel70_Valid_Out & channel57_Kernel70_Valid_Out & channel58_Kernel70_Valid_Out & channel59_Kernel70_Valid_Out & channel60_Kernel70_Valid_Out & channel61_Kernel70_Valid_Out & channel62_Kernel70_Valid_Out & channel63_Kernel70_Valid_Out & channel64_Kernel70_Valid_Out;

	wire channel1_Kernel71_Valid_Out, channel2_Kernel71_Valid_Out, channel3_Kernel71_Valid_Out, channel4_Kernel71_Valid_Out, channel5_Kernel71_Valid_Out, channel6_Kernel71_Valid_Out, channel7_Kernel71_Valid_Out, channel8_Kernel71_Valid_Out, channel9_Kernel71_Valid_Out, channel10_Kernel71_Valid_Out, channel11_Kernel71_Valid_Out, channel12_Kernel71_Valid_Out, channel13_Kernel71_Valid_Out, channel14_Kernel71_Valid_Out, channel15_Kernel71_Valid_Out, channel16_Kernel71_Valid_Out, channel17_Kernel71_Valid_Out, channel18_Kernel71_Valid_Out, channel19_Kernel71_Valid_Out, channel20_Kernel71_Valid_Out, channel21_Kernel71_Valid_Out, channel22_Kernel71_Valid_Out, channel23_Kernel71_Valid_Out, channel24_Kernel71_Valid_Out, channel25_Kernel71_Valid_Out, channel26_Kernel71_Valid_Out, channel27_Kernel71_Valid_Out, channel28_Kernel71_Valid_Out, channel29_Kernel71_Valid_Out, channel30_Kernel71_Valid_Out, channel31_Kernel71_Valid_Out, channel32_Kernel71_Valid_Out, channel33_Kernel71_Valid_Out, channel34_Kernel71_Valid_Out, channel35_Kernel71_Valid_Out, channel36_Kernel71_Valid_Out, channel37_Kernel71_Valid_Out, channel38_Kernel71_Valid_Out, channel39_Kernel71_Valid_Out, channel40_Kernel71_Valid_Out, channel41_Kernel71_Valid_Out, channel42_Kernel71_Valid_Out, channel43_Kernel71_Valid_Out, channel44_Kernel71_Valid_Out, channel45_Kernel71_Valid_Out, channel46_Kernel71_Valid_Out, channel47_Kernel71_Valid_Out, channel48_Kernel71_Valid_Out, channel49_Kernel71_Valid_Out, channel50_Kernel71_Valid_Out, channel51_Kernel71_Valid_Out, channel52_Kernel71_Valid_Out, channel53_Kernel71_Valid_Out, channel54_Kernel71_Valid_Out, channel55_Kernel71_Valid_Out, channel56_Kernel71_Valid_Out, channel57_Kernel71_Valid_Out, channel58_Kernel71_Valid_Out, channel59_Kernel71_Valid_Out, channel60_Kernel71_Valid_Out, channel61_Kernel71_Valid_Out, channel62_Kernel71_Valid_Out, channel63_Kernel71_Valid_Out, channel64_Kernel71_Valid_Out;

	assign add_kernel71=channel1_Kernel71_Valid_Out & channel2_Kernel71_Valid_Out & channel3_Kernel71_Valid_Out & channel4_Kernel71_Valid_Out & channel5_Kernel71_Valid_Out & channel6_Kernel71_Valid_Out & channel7_Kernel71_Valid_Out & channel8_Kernel71_Valid_Out & channel9_Kernel71_Valid_Out & channel10_Kernel71_Valid_Out & channel11_Kernel71_Valid_Out & channel12_Kernel71_Valid_Out & channel13_Kernel71_Valid_Out & channel14_Kernel71_Valid_Out & channel15_Kernel71_Valid_Out & channel16_Kernel71_Valid_Out & channel17_Kernel71_Valid_Out & channel18_Kernel71_Valid_Out & channel19_Kernel71_Valid_Out & channel20_Kernel71_Valid_Out & channel21_Kernel71_Valid_Out & channel22_Kernel71_Valid_Out & channel23_Kernel71_Valid_Out & channel24_Kernel71_Valid_Out & channel25_Kernel71_Valid_Out & channel26_Kernel71_Valid_Out & channel27_Kernel71_Valid_Out & channel28_Kernel71_Valid_Out & channel29_Kernel71_Valid_Out & channel30_Kernel71_Valid_Out & channel31_Kernel71_Valid_Out & channel32_Kernel71_Valid_Out & channel33_Kernel71_Valid_Out & channel34_Kernel71_Valid_Out & channel35_Kernel71_Valid_Out & channel36_Kernel71_Valid_Out & channel37_Kernel71_Valid_Out & channel38_Kernel71_Valid_Out & channel39_Kernel71_Valid_Out & channel40_Kernel71_Valid_Out & channel41_Kernel71_Valid_Out & channel42_Kernel71_Valid_Out & channel43_Kernel71_Valid_Out & channel44_Kernel71_Valid_Out & channel45_Kernel71_Valid_Out & channel46_Kernel71_Valid_Out & channel47_Kernel71_Valid_Out & channel48_Kernel71_Valid_Out & channel49_Kernel71_Valid_Out & channel50_Kernel71_Valid_Out & channel51_Kernel71_Valid_Out & channel52_Kernel71_Valid_Out & channel53_Kernel71_Valid_Out & channel54_Kernel71_Valid_Out & channel55_Kernel71_Valid_Out & channel56_Kernel71_Valid_Out & channel57_Kernel71_Valid_Out & channel58_Kernel71_Valid_Out & channel59_Kernel71_Valid_Out & channel60_Kernel71_Valid_Out & channel61_Kernel71_Valid_Out & channel62_Kernel71_Valid_Out & channel63_Kernel71_Valid_Out & channel64_Kernel71_Valid_Out;

	wire channel1_Kernel72_Valid_Out, channel2_Kernel72_Valid_Out, channel3_Kernel72_Valid_Out, channel4_Kernel72_Valid_Out, channel5_Kernel72_Valid_Out, channel6_Kernel72_Valid_Out, channel7_Kernel72_Valid_Out, channel8_Kernel72_Valid_Out, channel9_Kernel72_Valid_Out, channel10_Kernel72_Valid_Out, channel11_Kernel72_Valid_Out, channel12_Kernel72_Valid_Out, channel13_Kernel72_Valid_Out, channel14_Kernel72_Valid_Out, channel15_Kernel72_Valid_Out, channel16_Kernel72_Valid_Out, channel17_Kernel72_Valid_Out, channel18_Kernel72_Valid_Out, channel19_Kernel72_Valid_Out, channel20_Kernel72_Valid_Out, channel21_Kernel72_Valid_Out, channel22_Kernel72_Valid_Out, channel23_Kernel72_Valid_Out, channel24_Kernel72_Valid_Out, channel25_Kernel72_Valid_Out, channel26_Kernel72_Valid_Out, channel27_Kernel72_Valid_Out, channel28_Kernel72_Valid_Out, channel29_Kernel72_Valid_Out, channel30_Kernel72_Valid_Out, channel31_Kernel72_Valid_Out, channel32_Kernel72_Valid_Out, channel33_Kernel72_Valid_Out, channel34_Kernel72_Valid_Out, channel35_Kernel72_Valid_Out, channel36_Kernel72_Valid_Out, channel37_Kernel72_Valid_Out, channel38_Kernel72_Valid_Out, channel39_Kernel72_Valid_Out, channel40_Kernel72_Valid_Out, channel41_Kernel72_Valid_Out, channel42_Kernel72_Valid_Out, channel43_Kernel72_Valid_Out, channel44_Kernel72_Valid_Out, channel45_Kernel72_Valid_Out, channel46_Kernel72_Valid_Out, channel47_Kernel72_Valid_Out, channel48_Kernel72_Valid_Out, channel49_Kernel72_Valid_Out, channel50_Kernel72_Valid_Out, channel51_Kernel72_Valid_Out, channel52_Kernel72_Valid_Out, channel53_Kernel72_Valid_Out, channel54_Kernel72_Valid_Out, channel55_Kernel72_Valid_Out, channel56_Kernel72_Valid_Out, channel57_Kernel72_Valid_Out, channel58_Kernel72_Valid_Out, channel59_Kernel72_Valid_Out, channel60_Kernel72_Valid_Out, channel61_Kernel72_Valid_Out, channel62_Kernel72_Valid_Out, channel63_Kernel72_Valid_Out, channel64_Kernel72_Valid_Out;

	assign add_kernel72=channel1_Kernel72_Valid_Out & channel2_Kernel72_Valid_Out & channel3_Kernel72_Valid_Out & channel4_Kernel72_Valid_Out & channel5_Kernel72_Valid_Out & channel6_Kernel72_Valid_Out & channel7_Kernel72_Valid_Out & channel8_Kernel72_Valid_Out & channel9_Kernel72_Valid_Out & channel10_Kernel72_Valid_Out & channel11_Kernel72_Valid_Out & channel12_Kernel72_Valid_Out & channel13_Kernel72_Valid_Out & channel14_Kernel72_Valid_Out & channel15_Kernel72_Valid_Out & channel16_Kernel72_Valid_Out & channel17_Kernel72_Valid_Out & channel18_Kernel72_Valid_Out & channel19_Kernel72_Valid_Out & channel20_Kernel72_Valid_Out & channel21_Kernel72_Valid_Out & channel22_Kernel72_Valid_Out & channel23_Kernel72_Valid_Out & channel24_Kernel72_Valid_Out & channel25_Kernel72_Valid_Out & channel26_Kernel72_Valid_Out & channel27_Kernel72_Valid_Out & channel28_Kernel72_Valid_Out & channel29_Kernel72_Valid_Out & channel30_Kernel72_Valid_Out & channel31_Kernel72_Valid_Out & channel32_Kernel72_Valid_Out & channel33_Kernel72_Valid_Out & channel34_Kernel72_Valid_Out & channel35_Kernel72_Valid_Out & channel36_Kernel72_Valid_Out & channel37_Kernel72_Valid_Out & channel38_Kernel72_Valid_Out & channel39_Kernel72_Valid_Out & channel40_Kernel72_Valid_Out & channel41_Kernel72_Valid_Out & channel42_Kernel72_Valid_Out & channel43_Kernel72_Valid_Out & channel44_Kernel72_Valid_Out & channel45_Kernel72_Valid_Out & channel46_Kernel72_Valid_Out & channel47_Kernel72_Valid_Out & channel48_Kernel72_Valid_Out & channel49_Kernel72_Valid_Out & channel50_Kernel72_Valid_Out & channel51_Kernel72_Valid_Out & channel52_Kernel72_Valid_Out & channel53_Kernel72_Valid_Out & channel54_Kernel72_Valid_Out & channel55_Kernel72_Valid_Out & channel56_Kernel72_Valid_Out & channel57_Kernel72_Valid_Out & channel58_Kernel72_Valid_Out & channel59_Kernel72_Valid_Out & channel60_Kernel72_Valid_Out & channel61_Kernel72_Valid_Out & channel62_Kernel72_Valid_Out & channel63_Kernel72_Valid_Out & channel64_Kernel72_Valid_Out;

	wire channel1_Kernel73_Valid_Out, channel2_Kernel73_Valid_Out, channel3_Kernel73_Valid_Out, channel4_Kernel73_Valid_Out, channel5_Kernel73_Valid_Out, channel6_Kernel73_Valid_Out, channel7_Kernel73_Valid_Out, channel8_Kernel73_Valid_Out, channel9_Kernel73_Valid_Out, channel10_Kernel73_Valid_Out, channel11_Kernel73_Valid_Out, channel12_Kernel73_Valid_Out, channel13_Kernel73_Valid_Out, channel14_Kernel73_Valid_Out, channel15_Kernel73_Valid_Out, channel16_Kernel73_Valid_Out, channel17_Kernel73_Valid_Out, channel18_Kernel73_Valid_Out, channel19_Kernel73_Valid_Out, channel20_Kernel73_Valid_Out, channel21_Kernel73_Valid_Out, channel22_Kernel73_Valid_Out, channel23_Kernel73_Valid_Out, channel24_Kernel73_Valid_Out, channel25_Kernel73_Valid_Out, channel26_Kernel73_Valid_Out, channel27_Kernel73_Valid_Out, channel28_Kernel73_Valid_Out, channel29_Kernel73_Valid_Out, channel30_Kernel73_Valid_Out, channel31_Kernel73_Valid_Out, channel32_Kernel73_Valid_Out, channel33_Kernel73_Valid_Out, channel34_Kernel73_Valid_Out, channel35_Kernel73_Valid_Out, channel36_Kernel73_Valid_Out, channel37_Kernel73_Valid_Out, channel38_Kernel73_Valid_Out, channel39_Kernel73_Valid_Out, channel40_Kernel73_Valid_Out, channel41_Kernel73_Valid_Out, channel42_Kernel73_Valid_Out, channel43_Kernel73_Valid_Out, channel44_Kernel73_Valid_Out, channel45_Kernel73_Valid_Out, channel46_Kernel73_Valid_Out, channel47_Kernel73_Valid_Out, channel48_Kernel73_Valid_Out, channel49_Kernel73_Valid_Out, channel50_Kernel73_Valid_Out, channel51_Kernel73_Valid_Out, channel52_Kernel73_Valid_Out, channel53_Kernel73_Valid_Out, channel54_Kernel73_Valid_Out, channel55_Kernel73_Valid_Out, channel56_Kernel73_Valid_Out, channel57_Kernel73_Valid_Out, channel58_Kernel73_Valid_Out, channel59_Kernel73_Valid_Out, channel60_Kernel73_Valid_Out, channel61_Kernel73_Valid_Out, channel62_Kernel73_Valid_Out, channel63_Kernel73_Valid_Out, channel64_Kernel73_Valid_Out;

	assign add_kernel73=channel1_Kernel73_Valid_Out & channel2_Kernel73_Valid_Out & channel3_Kernel73_Valid_Out & channel4_Kernel73_Valid_Out & channel5_Kernel73_Valid_Out & channel6_Kernel73_Valid_Out & channel7_Kernel73_Valid_Out & channel8_Kernel73_Valid_Out & channel9_Kernel73_Valid_Out & channel10_Kernel73_Valid_Out & channel11_Kernel73_Valid_Out & channel12_Kernel73_Valid_Out & channel13_Kernel73_Valid_Out & channel14_Kernel73_Valid_Out & channel15_Kernel73_Valid_Out & channel16_Kernel73_Valid_Out & channel17_Kernel73_Valid_Out & channel18_Kernel73_Valid_Out & channel19_Kernel73_Valid_Out & channel20_Kernel73_Valid_Out & channel21_Kernel73_Valid_Out & channel22_Kernel73_Valid_Out & channel23_Kernel73_Valid_Out & channel24_Kernel73_Valid_Out & channel25_Kernel73_Valid_Out & channel26_Kernel73_Valid_Out & channel27_Kernel73_Valid_Out & channel28_Kernel73_Valid_Out & channel29_Kernel73_Valid_Out & channel30_Kernel73_Valid_Out & channel31_Kernel73_Valid_Out & channel32_Kernel73_Valid_Out & channel33_Kernel73_Valid_Out & channel34_Kernel73_Valid_Out & channel35_Kernel73_Valid_Out & channel36_Kernel73_Valid_Out & channel37_Kernel73_Valid_Out & channel38_Kernel73_Valid_Out & channel39_Kernel73_Valid_Out & channel40_Kernel73_Valid_Out & channel41_Kernel73_Valid_Out & channel42_Kernel73_Valid_Out & channel43_Kernel73_Valid_Out & channel44_Kernel73_Valid_Out & channel45_Kernel73_Valid_Out & channel46_Kernel73_Valid_Out & channel47_Kernel73_Valid_Out & channel48_Kernel73_Valid_Out & channel49_Kernel73_Valid_Out & channel50_Kernel73_Valid_Out & channel51_Kernel73_Valid_Out & channel52_Kernel73_Valid_Out & channel53_Kernel73_Valid_Out & channel54_Kernel73_Valid_Out & channel55_Kernel73_Valid_Out & channel56_Kernel73_Valid_Out & channel57_Kernel73_Valid_Out & channel58_Kernel73_Valid_Out & channel59_Kernel73_Valid_Out & channel60_Kernel73_Valid_Out & channel61_Kernel73_Valid_Out & channel62_Kernel73_Valid_Out & channel63_Kernel73_Valid_Out & channel64_Kernel73_Valid_Out;

	wire channel1_Kernel74_Valid_Out, channel2_Kernel74_Valid_Out, channel3_Kernel74_Valid_Out, channel4_Kernel74_Valid_Out, channel5_Kernel74_Valid_Out, channel6_Kernel74_Valid_Out, channel7_Kernel74_Valid_Out, channel8_Kernel74_Valid_Out, channel9_Kernel74_Valid_Out, channel10_Kernel74_Valid_Out, channel11_Kernel74_Valid_Out, channel12_Kernel74_Valid_Out, channel13_Kernel74_Valid_Out, channel14_Kernel74_Valid_Out, channel15_Kernel74_Valid_Out, channel16_Kernel74_Valid_Out, channel17_Kernel74_Valid_Out, channel18_Kernel74_Valid_Out, channel19_Kernel74_Valid_Out, channel20_Kernel74_Valid_Out, channel21_Kernel74_Valid_Out, channel22_Kernel74_Valid_Out, channel23_Kernel74_Valid_Out, channel24_Kernel74_Valid_Out, channel25_Kernel74_Valid_Out, channel26_Kernel74_Valid_Out, channel27_Kernel74_Valid_Out, channel28_Kernel74_Valid_Out, channel29_Kernel74_Valid_Out, channel30_Kernel74_Valid_Out, channel31_Kernel74_Valid_Out, channel32_Kernel74_Valid_Out, channel33_Kernel74_Valid_Out, channel34_Kernel74_Valid_Out, channel35_Kernel74_Valid_Out, channel36_Kernel74_Valid_Out, channel37_Kernel74_Valid_Out, channel38_Kernel74_Valid_Out, channel39_Kernel74_Valid_Out, channel40_Kernel74_Valid_Out, channel41_Kernel74_Valid_Out, channel42_Kernel74_Valid_Out, channel43_Kernel74_Valid_Out, channel44_Kernel74_Valid_Out, channel45_Kernel74_Valid_Out, channel46_Kernel74_Valid_Out, channel47_Kernel74_Valid_Out, channel48_Kernel74_Valid_Out, channel49_Kernel74_Valid_Out, channel50_Kernel74_Valid_Out, channel51_Kernel74_Valid_Out, channel52_Kernel74_Valid_Out, channel53_Kernel74_Valid_Out, channel54_Kernel74_Valid_Out, channel55_Kernel74_Valid_Out, channel56_Kernel74_Valid_Out, channel57_Kernel74_Valid_Out, channel58_Kernel74_Valid_Out, channel59_Kernel74_Valid_Out, channel60_Kernel74_Valid_Out, channel61_Kernel74_Valid_Out, channel62_Kernel74_Valid_Out, channel63_Kernel74_Valid_Out, channel64_Kernel74_Valid_Out;

	assign add_kernel74=channel1_Kernel74_Valid_Out & channel2_Kernel74_Valid_Out & channel3_Kernel74_Valid_Out & channel4_Kernel74_Valid_Out & channel5_Kernel74_Valid_Out & channel6_Kernel74_Valid_Out & channel7_Kernel74_Valid_Out & channel8_Kernel74_Valid_Out & channel9_Kernel74_Valid_Out & channel10_Kernel74_Valid_Out & channel11_Kernel74_Valid_Out & channel12_Kernel74_Valid_Out & channel13_Kernel74_Valid_Out & channel14_Kernel74_Valid_Out & channel15_Kernel74_Valid_Out & channel16_Kernel74_Valid_Out & channel17_Kernel74_Valid_Out & channel18_Kernel74_Valid_Out & channel19_Kernel74_Valid_Out & channel20_Kernel74_Valid_Out & channel21_Kernel74_Valid_Out & channel22_Kernel74_Valid_Out & channel23_Kernel74_Valid_Out & channel24_Kernel74_Valid_Out & channel25_Kernel74_Valid_Out & channel26_Kernel74_Valid_Out & channel27_Kernel74_Valid_Out & channel28_Kernel74_Valid_Out & channel29_Kernel74_Valid_Out & channel30_Kernel74_Valid_Out & channel31_Kernel74_Valid_Out & channel32_Kernel74_Valid_Out & channel33_Kernel74_Valid_Out & channel34_Kernel74_Valid_Out & channel35_Kernel74_Valid_Out & channel36_Kernel74_Valid_Out & channel37_Kernel74_Valid_Out & channel38_Kernel74_Valid_Out & channel39_Kernel74_Valid_Out & channel40_Kernel74_Valid_Out & channel41_Kernel74_Valid_Out & channel42_Kernel74_Valid_Out & channel43_Kernel74_Valid_Out & channel44_Kernel74_Valid_Out & channel45_Kernel74_Valid_Out & channel46_Kernel74_Valid_Out & channel47_Kernel74_Valid_Out & channel48_Kernel74_Valid_Out & channel49_Kernel74_Valid_Out & channel50_Kernel74_Valid_Out & channel51_Kernel74_Valid_Out & channel52_Kernel74_Valid_Out & channel53_Kernel74_Valid_Out & channel54_Kernel74_Valid_Out & channel55_Kernel74_Valid_Out & channel56_Kernel74_Valid_Out & channel57_Kernel74_Valid_Out & channel58_Kernel74_Valid_Out & channel59_Kernel74_Valid_Out & channel60_Kernel74_Valid_Out & channel61_Kernel74_Valid_Out & channel62_Kernel74_Valid_Out & channel63_Kernel74_Valid_Out & channel64_Kernel74_Valid_Out;

	wire channel1_Kernel75_Valid_Out, channel2_Kernel75_Valid_Out, channel3_Kernel75_Valid_Out, channel4_Kernel75_Valid_Out, channel5_Kernel75_Valid_Out, channel6_Kernel75_Valid_Out, channel7_Kernel75_Valid_Out, channel8_Kernel75_Valid_Out, channel9_Kernel75_Valid_Out, channel10_Kernel75_Valid_Out, channel11_Kernel75_Valid_Out, channel12_Kernel75_Valid_Out, channel13_Kernel75_Valid_Out, channel14_Kernel75_Valid_Out, channel15_Kernel75_Valid_Out, channel16_Kernel75_Valid_Out, channel17_Kernel75_Valid_Out, channel18_Kernel75_Valid_Out, channel19_Kernel75_Valid_Out, channel20_Kernel75_Valid_Out, channel21_Kernel75_Valid_Out, channel22_Kernel75_Valid_Out, channel23_Kernel75_Valid_Out, channel24_Kernel75_Valid_Out, channel25_Kernel75_Valid_Out, channel26_Kernel75_Valid_Out, channel27_Kernel75_Valid_Out, channel28_Kernel75_Valid_Out, channel29_Kernel75_Valid_Out, channel30_Kernel75_Valid_Out, channel31_Kernel75_Valid_Out, channel32_Kernel75_Valid_Out, channel33_Kernel75_Valid_Out, channel34_Kernel75_Valid_Out, channel35_Kernel75_Valid_Out, channel36_Kernel75_Valid_Out, channel37_Kernel75_Valid_Out, channel38_Kernel75_Valid_Out, channel39_Kernel75_Valid_Out, channel40_Kernel75_Valid_Out, channel41_Kernel75_Valid_Out, channel42_Kernel75_Valid_Out, channel43_Kernel75_Valid_Out, channel44_Kernel75_Valid_Out, channel45_Kernel75_Valid_Out, channel46_Kernel75_Valid_Out, channel47_Kernel75_Valid_Out, channel48_Kernel75_Valid_Out, channel49_Kernel75_Valid_Out, channel50_Kernel75_Valid_Out, channel51_Kernel75_Valid_Out, channel52_Kernel75_Valid_Out, channel53_Kernel75_Valid_Out, channel54_Kernel75_Valid_Out, channel55_Kernel75_Valid_Out, channel56_Kernel75_Valid_Out, channel57_Kernel75_Valid_Out, channel58_Kernel75_Valid_Out, channel59_Kernel75_Valid_Out, channel60_Kernel75_Valid_Out, channel61_Kernel75_Valid_Out, channel62_Kernel75_Valid_Out, channel63_Kernel75_Valid_Out, channel64_Kernel75_Valid_Out;

	assign add_kernel75=channel1_Kernel75_Valid_Out & channel2_Kernel75_Valid_Out & channel3_Kernel75_Valid_Out & channel4_Kernel75_Valid_Out & channel5_Kernel75_Valid_Out & channel6_Kernel75_Valid_Out & channel7_Kernel75_Valid_Out & channel8_Kernel75_Valid_Out & channel9_Kernel75_Valid_Out & channel10_Kernel75_Valid_Out & channel11_Kernel75_Valid_Out & channel12_Kernel75_Valid_Out & channel13_Kernel75_Valid_Out & channel14_Kernel75_Valid_Out & channel15_Kernel75_Valid_Out & channel16_Kernel75_Valid_Out & channel17_Kernel75_Valid_Out & channel18_Kernel75_Valid_Out & channel19_Kernel75_Valid_Out & channel20_Kernel75_Valid_Out & channel21_Kernel75_Valid_Out & channel22_Kernel75_Valid_Out & channel23_Kernel75_Valid_Out & channel24_Kernel75_Valid_Out & channel25_Kernel75_Valid_Out & channel26_Kernel75_Valid_Out & channel27_Kernel75_Valid_Out & channel28_Kernel75_Valid_Out & channel29_Kernel75_Valid_Out & channel30_Kernel75_Valid_Out & channel31_Kernel75_Valid_Out & channel32_Kernel75_Valid_Out & channel33_Kernel75_Valid_Out & channel34_Kernel75_Valid_Out & channel35_Kernel75_Valid_Out & channel36_Kernel75_Valid_Out & channel37_Kernel75_Valid_Out & channel38_Kernel75_Valid_Out & channel39_Kernel75_Valid_Out & channel40_Kernel75_Valid_Out & channel41_Kernel75_Valid_Out & channel42_Kernel75_Valid_Out & channel43_Kernel75_Valid_Out & channel44_Kernel75_Valid_Out & channel45_Kernel75_Valid_Out & channel46_Kernel75_Valid_Out & channel47_Kernel75_Valid_Out & channel48_Kernel75_Valid_Out & channel49_Kernel75_Valid_Out & channel50_Kernel75_Valid_Out & channel51_Kernel75_Valid_Out & channel52_Kernel75_Valid_Out & channel53_Kernel75_Valid_Out & channel54_Kernel75_Valid_Out & channel55_Kernel75_Valid_Out & channel56_Kernel75_Valid_Out & channel57_Kernel75_Valid_Out & channel58_Kernel75_Valid_Out & channel59_Kernel75_Valid_Out & channel60_Kernel75_Valid_Out & channel61_Kernel75_Valid_Out & channel62_Kernel75_Valid_Out & channel63_Kernel75_Valid_Out & channel64_Kernel75_Valid_Out;

	wire channel1_Kernel76_Valid_Out, channel2_Kernel76_Valid_Out, channel3_Kernel76_Valid_Out, channel4_Kernel76_Valid_Out, channel5_Kernel76_Valid_Out, channel6_Kernel76_Valid_Out, channel7_Kernel76_Valid_Out, channel8_Kernel76_Valid_Out, channel9_Kernel76_Valid_Out, channel10_Kernel76_Valid_Out, channel11_Kernel76_Valid_Out, channel12_Kernel76_Valid_Out, channel13_Kernel76_Valid_Out, channel14_Kernel76_Valid_Out, channel15_Kernel76_Valid_Out, channel16_Kernel76_Valid_Out, channel17_Kernel76_Valid_Out, channel18_Kernel76_Valid_Out, channel19_Kernel76_Valid_Out, channel20_Kernel76_Valid_Out, channel21_Kernel76_Valid_Out, channel22_Kernel76_Valid_Out, channel23_Kernel76_Valid_Out, channel24_Kernel76_Valid_Out, channel25_Kernel76_Valid_Out, channel26_Kernel76_Valid_Out, channel27_Kernel76_Valid_Out, channel28_Kernel76_Valid_Out, channel29_Kernel76_Valid_Out, channel30_Kernel76_Valid_Out, channel31_Kernel76_Valid_Out, channel32_Kernel76_Valid_Out, channel33_Kernel76_Valid_Out, channel34_Kernel76_Valid_Out, channel35_Kernel76_Valid_Out, channel36_Kernel76_Valid_Out, channel37_Kernel76_Valid_Out, channel38_Kernel76_Valid_Out, channel39_Kernel76_Valid_Out, channel40_Kernel76_Valid_Out, channel41_Kernel76_Valid_Out, channel42_Kernel76_Valid_Out, channel43_Kernel76_Valid_Out, channel44_Kernel76_Valid_Out, channel45_Kernel76_Valid_Out, channel46_Kernel76_Valid_Out, channel47_Kernel76_Valid_Out, channel48_Kernel76_Valid_Out, channel49_Kernel76_Valid_Out, channel50_Kernel76_Valid_Out, channel51_Kernel76_Valid_Out, channel52_Kernel76_Valid_Out, channel53_Kernel76_Valid_Out, channel54_Kernel76_Valid_Out, channel55_Kernel76_Valid_Out, channel56_Kernel76_Valid_Out, channel57_Kernel76_Valid_Out, channel58_Kernel76_Valid_Out, channel59_Kernel76_Valid_Out, channel60_Kernel76_Valid_Out, channel61_Kernel76_Valid_Out, channel62_Kernel76_Valid_Out, channel63_Kernel76_Valid_Out, channel64_Kernel76_Valid_Out;

	assign add_kernel76=channel1_Kernel76_Valid_Out & channel2_Kernel76_Valid_Out & channel3_Kernel76_Valid_Out & channel4_Kernel76_Valid_Out & channel5_Kernel76_Valid_Out & channel6_Kernel76_Valid_Out & channel7_Kernel76_Valid_Out & channel8_Kernel76_Valid_Out & channel9_Kernel76_Valid_Out & channel10_Kernel76_Valid_Out & channel11_Kernel76_Valid_Out & channel12_Kernel76_Valid_Out & channel13_Kernel76_Valid_Out & channel14_Kernel76_Valid_Out & channel15_Kernel76_Valid_Out & channel16_Kernel76_Valid_Out & channel17_Kernel76_Valid_Out & channel18_Kernel76_Valid_Out & channel19_Kernel76_Valid_Out & channel20_Kernel76_Valid_Out & channel21_Kernel76_Valid_Out & channel22_Kernel76_Valid_Out & channel23_Kernel76_Valid_Out & channel24_Kernel76_Valid_Out & channel25_Kernel76_Valid_Out & channel26_Kernel76_Valid_Out & channel27_Kernel76_Valid_Out & channel28_Kernel76_Valid_Out & channel29_Kernel76_Valid_Out & channel30_Kernel76_Valid_Out & channel31_Kernel76_Valid_Out & channel32_Kernel76_Valid_Out & channel33_Kernel76_Valid_Out & channel34_Kernel76_Valid_Out & channel35_Kernel76_Valid_Out & channel36_Kernel76_Valid_Out & channel37_Kernel76_Valid_Out & channel38_Kernel76_Valid_Out & channel39_Kernel76_Valid_Out & channel40_Kernel76_Valid_Out & channel41_Kernel76_Valid_Out & channel42_Kernel76_Valid_Out & channel43_Kernel76_Valid_Out & channel44_Kernel76_Valid_Out & channel45_Kernel76_Valid_Out & channel46_Kernel76_Valid_Out & channel47_Kernel76_Valid_Out & channel48_Kernel76_Valid_Out & channel49_Kernel76_Valid_Out & channel50_Kernel76_Valid_Out & channel51_Kernel76_Valid_Out & channel52_Kernel76_Valid_Out & channel53_Kernel76_Valid_Out & channel54_Kernel76_Valid_Out & channel55_Kernel76_Valid_Out & channel56_Kernel76_Valid_Out & channel57_Kernel76_Valid_Out & channel58_Kernel76_Valid_Out & channel59_Kernel76_Valid_Out & channel60_Kernel76_Valid_Out & channel61_Kernel76_Valid_Out & channel62_Kernel76_Valid_Out & channel63_Kernel76_Valid_Out & channel64_Kernel76_Valid_Out;

	wire channel1_Kernel77_Valid_Out, channel2_Kernel77_Valid_Out, channel3_Kernel77_Valid_Out, channel4_Kernel77_Valid_Out, channel5_Kernel77_Valid_Out, channel6_Kernel77_Valid_Out, channel7_Kernel77_Valid_Out, channel8_Kernel77_Valid_Out, channel9_Kernel77_Valid_Out, channel10_Kernel77_Valid_Out, channel11_Kernel77_Valid_Out, channel12_Kernel77_Valid_Out, channel13_Kernel77_Valid_Out, channel14_Kernel77_Valid_Out, channel15_Kernel77_Valid_Out, channel16_Kernel77_Valid_Out, channel17_Kernel77_Valid_Out, channel18_Kernel77_Valid_Out, channel19_Kernel77_Valid_Out, channel20_Kernel77_Valid_Out, channel21_Kernel77_Valid_Out, channel22_Kernel77_Valid_Out, channel23_Kernel77_Valid_Out, channel24_Kernel77_Valid_Out, channel25_Kernel77_Valid_Out, channel26_Kernel77_Valid_Out, channel27_Kernel77_Valid_Out, channel28_Kernel77_Valid_Out, channel29_Kernel77_Valid_Out, channel30_Kernel77_Valid_Out, channel31_Kernel77_Valid_Out, channel32_Kernel77_Valid_Out, channel33_Kernel77_Valid_Out, channel34_Kernel77_Valid_Out, channel35_Kernel77_Valid_Out, channel36_Kernel77_Valid_Out, channel37_Kernel77_Valid_Out, channel38_Kernel77_Valid_Out, channel39_Kernel77_Valid_Out, channel40_Kernel77_Valid_Out, channel41_Kernel77_Valid_Out, channel42_Kernel77_Valid_Out, channel43_Kernel77_Valid_Out, channel44_Kernel77_Valid_Out, channel45_Kernel77_Valid_Out, channel46_Kernel77_Valid_Out, channel47_Kernel77_Valid_Out, channel48_Kernel77_Valid_Out, channel49_Kernel77_Valid_Out, channel50_Kernel77_Valid_Out, channel51_Kernel77_Valid_Out, channel52_Kernel77_Valid_Out, channel53_Kernel77_Valid_Out, channel54_Kernel77_Valid_Out, channel55_Kernel77_Valid_Out, channel56_Kernel77_Valid_Out, channel57_Kernel77_Valid_Out, channel58_Kernel77_Valid_Out, channel59_Kernel77_Valid_Out, channel60_Kernel77_Valid_Out, channel61_Kernel77_Valid_Out, channel62_Kernel77_Valid_Out, channel63_Kernel77_Valid_Out, channel64_Kernel77_Valid_Out;

	assign add_kernel77=channel1_Kernel77_Valid_Out & channel2_Kernel77_Valid_Out & channel3_Kernel77_Valid_Out & channel4_Kernel77_Valid_Out & channel5_Kernel77_Valid_Out & channel6_Kernel77_Valid_Out & channel7_Kernel77_Valid_Out & channel8_Kernel77_Valid_Out & channel9_Kernel77_Valid_Out & channel10_Kernel77_Valid_Out & channel11_Kernel77_Valid_Out & channel12_Kernel77_Valid_Out & channel13_Kernel77_Valid_Out & channel14_Kernel77_Valid_Out & channel15_Kernel77_Valid_Out & channel16_Kernel77_Valid_Out & channel17_Kernel77_Valid_Out & channel18_Kernel77_Valid_Out & channel19_Kernel77_Valid_Out & channel20_Kernel77_Valid_Out & channel21_Kernel77_Valid_Out & channel22_Kernel77_Valid_Out & channel23_Kernel77_Valid_Out & channel24_Kernel77_Valid_Out & channel25_Kernel77_Valid_Out & channel26_Kernel77_Valid_Out & channel27_Kernel77_Valid_Out & channel28_Kernel77_Valid_Out & channel29_Kernel77_Valid_Out & channel30_Kernel77_Valid_Out & channel31_Kernel77_Valid_Out & channel32_Kernel77_Valid_Out & channel33_Kernel77_Valid_Out & channel34_Kernel77_Valid_Out & channel35_Kernel77_Valid_Out & channel36_Kernel77_Valid_Out & channel37_Kernel77_Valid_Out & channel38_Kernel77_Valid_Out & channel39_Kernel77_Valid_Out & channel40_Kernel77_Valid_Out & channel41_Kernel77_Valid_Out & channel42_Kernel77_Valid_Out & channel43_Kernel77_Valid_Out & channel44_Kernel77_Valid_Out & channel45_Kernel77_Valid_Out & channel46_Kernel77_Valid_Out & channel47_Kernel77_Valid_Out & channel48_Kernel77_Valid_Out & channel49_Kernel77_Valid_Out & channel50_Kernel77_Valid_Out & channel51_Kernel77_Valid_Out & channel52_Kernel77_Valid_Out & channel53_Kernel77_Valid_Out & channel54_Kernel77_Valid_Out & channel55_Kernel77_Valid_Out & channel56_Kernel77_Valid_Out & channel57_Kernel77_Valid_Out & channel58_Kernel77_Valid_Out & channel59_Kernel77_Valid_Out & channel60_Kernel77_Valid_Out & channel61_Kernel77_Valid_Out & channel62_Kernel77_Valid_Out & channel63_Kernel77_Valid_Out & channel64_Kernel77_Valid_Out;

	wire channel1_Kernel78_Valid_Out, channel2_Kernel78_Valid_Out, channel3_Kernel78_Valid_Out, channel4_Kernel78_Valid_Out, channel5_Kernel78_Valid_Out, channel6_Kernel78_Valid_Out, channel7_Kernel78_Valid_Out, channel8_Kernel78_Valid_Out, channel9_Kernel78_Valid_Out, channel10_Kernel78_Valid_Out, channel11_Kernel78_Valid_Out, channel12_Kernel78_Valid_Out, channel13_Kernel78_Valid_Out, channel14_Kernel78_Valid_Out, channel15_Kernel78_Valid_Out, channel16_Kernel78_Valid_Out, channel17_Kernel78_Valid_Out, channel18_Kernel78_Valid_Out, channel19_Kernel78_Valid_Out, channel20_Kernel78_Valid_Out, channel21_Kernel78_Valid_Out, channel22_Kernel78_Valid_Out, channel23_Kernel78_Valid_Out, channel24_Kernel78_Valid_Out, channel25_Kernel78_Valid_Out, channel26_Kernel78_Valid_Out, channel27_Kernel78_Valid_Out, channel28_Kernel78_Valid_Out, channel29_Kernel78_Valid_Out, channel30_Kernel78_Valid_Out, channel31_Kernel78_Valid_Out, channel32_Kernel78_Valid_Out, channel33_Kernel78_Valid_Out, channel34_Kernel78_Valid_Out, channel35_Kernel78_Valid_Out, channel36_Kernel78_Valid_Out, channel37_Kernel78_Valid_Out, channel38_Kernel78_Valid_Out, channel39_Kernel78_Valid_Out, channel40_Kernel78_Valid_Out, channel41_Kernel78_Valid_Out, channel42_Kernel78_Valid_Out, channel43_Kernel78_Valid_Out, channel44_Kernel78_Valid_Out, channel45_Kernel78_Valid_Out, channel46_Kernel78_Valid_Out, channel47_Kernel78_Valid_Out, channel48_Kernel78_Valid_Out, channel49_Kernel78_Valid_Out, channel50_Kernel78_Valid_Out, channel51_Kernel78_Valid_Out, channel52_Kernel78_Valid_Out, channel53_Kernel78_Valid_Out, channel54_Kernel78_Valid_Out, channel55_Kernel78_Valid_Out, channel56_Kernel78_Valid_Out, channel57_Kernel78_Valid_Out, channel58_Kernel78_Valid_Out, channel59_Kernel78_Valid_Out, channel60_Kernel78_Valid_Out, channel61_Kernel78_Valid_Out, channel62_Kernel78_Valid_Out, channel63_Kernel78_Valid_Out, channel64_Kernel78_Valid_Out;

	assign add_kernel78=channel1_Kernel78_Valid_Out & channel2_Kernel78_Valid_Out & channel3_Kernel78_Valid_Out & channel4_Kernel78_Valid_Out & channel5_Kernel78_Valid_Out & channel6_Kernel78_Valid_Out & channel7_Kernel78_Valid_Out & channel8_Kernel78_Valid_Out & channel9_Kernel78_Valid_Out & channel10_Kernel78_Valid_Out & channel11_Kernel78_Valid_Out & channel12_Kernel78_Valid_Out & channel13_Kernel78_Valid_Out & channel14_Kernel78_Valid_Out & channel15_Kernel78_Valid_Out & channel16_Kernel78_Valid_Out & channel17_Kernel78_Valid_Out & channel18_Kernel78_Valid_Out & channel19_Kernel78_Valid_Out & channel20_Kernel78_Valid_Out & channel21_Kernel78_Valid_Out & channel22_Kernel78_Valid_Out & channel23_Kernel78_Valid_Out & channel24_Kernel78_Valid_Out & channel25_Kernel78_Valid_Out & channel26_Kernel78_Valid_Out & channel27_Kernel78_Valid_Out & channel28_Kernel78_Valid_Out & channel29_Kernel78_Valid_Out & channel30_Kernel78_Valid_Out & channel31_Kernel78_Valid_Out & channel32_Kernel78_Valid_Out & channel33_Kernel78_Valid_Out & channel34_Kernel78_Valid_Out & channel35_Kernel78_Valid_Out & channel36_Kernel78_Valid_Out & channel37_Kernel78_Valid_Out & channel38_Kernel78_Valid_Out & channel39_Kernel78_Valid_Out & channel40_Kernel78_Valid_Out & channel41_Kernel78_Valid_Out & channel42_Kernel78_Valid_Out & channel43_Kernel78_Valid_Out & channel44_Kernel78_Valid_Out & channel45_Kernel78_Valid_Out & channel46_Kernel78_Valid_Out & channel47_Kernel78_Valid_Out & channel48_Kernel78_Valid_Out & channel49_Kernel78_Valid_Out & channel50_Kernel78_Valid_Out & channel51_Kernel78_Valid_Out & channel52_Kernel78_Valid_Out & channel53_Kernel78_Valid_Out & channel54_Kernel78_Valid_Out & channel55_Kernel78_Valid_Out & channel56_Kernel78_Valid_Out & channel57_Kernel78_Valid_Out & channel58_Kernel78_Valid_Out & channel59_Kernel78_Valid_Out & channel60_Kernel78_Valid_Out & channel61_Kernel78_Valid_Out & channel62_Kernel78_Valid_Out & channel63_Kernel78_Valid_Out & channel64_Kernel78_Valid_Out;

	wire channel1_Kernel79_Valid_Out, channel2_Kernel79_Valid_Out, channel3_Kernel79_Valid_Out, channel4_Kernel79_Valid_Out, channel5_Kernel79_Valid_Out, channel6_Kernel79_Valid_Out, channel7_Kernel79_Valid_Out, channel8_Kernel79_Valid_Out, channel9_Kernel79_Valid_Out, channel10_Kernel79_Valid_Out, channel11_Kernel79_Valid_Out, channel12_Kernel79_Valid_Out, channel13_Kernel79_Valid_Out, channel14_Kernel79_Valid_Out, channel15_Kernel79_Valid_Out, channel16_Kernel79_Valid_Out, channel17_Kernel79_Valid_Out, channel18_Kernel79_Valid_Out, channel19_Kernel79_Valid_Out, channel20_Kernel79_Valid_Out, channel21_Kernel79_Valid_Out, channel22_Kernel79_Valid_Out, channel23_Kernel79_Valid_Out, channel24_Kernel79_Valid_Out, channel25_Kernel79_Valid_Out, channel26_Kernel79_Valid_Out, channel27_Kernel79_Valid_Out, channel28_Kernel79_Valid_Out, channel29_Kernel79_Valid_Out, channel30_Kernel79_Valid_Out, channel31_Kernel79_Valid_Out, channel32_Kernel79_Valid_Out, channel33_Kernel79_Valid_Out, channel34_Kernel79_Valid_Out, channel35_Kernel79_Valid_Out, channel36_Kernel79_Valid_Out, channel37_Kernel79_Valid_Out, channel38_Kernel79_Valid_Out, channel39_Kernel79_Valid_Out, channel40_Kernel79_Valid_Out, channel41_Kernel79_Valid_Out, channel42_Kernel79_Valid_Out, channel43_Kernel79_Valid_Out, channel44_Kernel79_Valid_Out, channel45_Kernel79_Valid_Out, channel46_Kernel79_Valid_Out, channel47_Kernel79_Valid_Out, channel48_Kernel79_Valid_Out, channel49_Kernel79_Valid_Out, channel50_Kernel79_Valid_Out, channel51_Kernel79_Valid_Out, channel52_Kernel79_Valid_Out, channel53_Kernel79_Valid_Out, channel54_Kernel79_Valid_Out, channel55_Kernel79_Valid_Out, channel56_Kernel79_Valid_Out, channel57_Kernel79_Valid_Out, channel58_Kernel79_Valid_Out, channel59_Kernel79_Valid_Out, channel60_Kernel79_Valid_Out, channel61_Kernel79_Valid_Out, channel62_Kernel79_Valid_Out, channel63_Kernel79_Valid_Out, channel64_Kernel79_Valid_Out;

	assign add_kernel79=channel1_Kernel79_Valid_Out & channel2_Kernel79_Valid_Out & channel3_Kernel79_Valid_Out & channel4_Kernel79_Valid_Out & channel5_Kernel79_Valid_Out & channel6_Kernel79_Valid_Out & channel7_Kernel79_Valid_Out & channel8_Kernel79_Valid_Out & channel9_Kernel79_Valid_Out & channel10_Kernel79_Valid_Out & channel11_Kernel79_Valid_Out & channel12_Kernel79_Valid_Out & channel13_Kernel79_Valid_Out & channel14_Kernel79_Valid_Out & channel15_Kernel79_Valid_Out & channel16_Kernel79_Valid_Out & channel17_Kernel79_Valid_Out & channel18_Kernel79_Valid_Out & channel19_Kernel79_Valid_Out & channel20_Kernel79_Valid_Out & channel21_Kernel79_Valid_Out & channel22_Kernel79_Valid_Out & channel23_Kernel79_Valid_Out & channel24_Kernel79_Valid_Out & channel25_Kernel79_Valid_Out & channel26_Kernel79_Valid_Out & channel27_Kernel79_Valid_Out & channel28_Kernel79_Valid_Out & channel29_Kernel79_Valid_Out & channel30_Kernel79_Valid_Out & channel31_Kernel79_Valid_Out & channel32_Kernel79_Valid_Out & channel33_Kernel79_Valid_Out & channel34_Kernel79_Valid_Out & channel35_Kernel79_Valid_Out & channel36_Kernel79_Valid_Out & channel37_Kernel79_Valid_Out & channel38_Kernel79_Valid_Out & channel39_Kernel79_Valid_Out & channel40_Kernel79_Valid_Out & channel41_Kernel79_Valid_Out & channel42_Kernel79_Valid_Out & channel43_Kernel79_Valid_Out & channel44_Kernel79_Valid_Out & channel45_Kernel79_Valid_Out & channel46_Kernel79_Valid_Out & channel47_Kernel79_Valid_Out & channel48_Kernel79_Valid_Out & channel49_Kernel79_Valid_Out & channel50_Kernel79_Valid_Out & channel51_Kernel79_Valid_Out & channel52_Kernel79_Valid_Out & channel53_Kernel79_Valid_Out & channel54_Kernel79_Valid_Out & channel55_Kernel79_Valid_Out & channel56_Kernel79_Valid_Out & channel57_Kernel79_Valid_Out & channel58_Kernel79_Valid_Out & channel59_Kernel79_Valid_Out & channel60_Kernel79_Valid_Out & channel61_Kernel79_Valid_Out & channel62_Kernel79_Valid_Out & channel63_Kernel79_Valid_Out & channel64_Kernel79_Valid_Out;

	wire channel1_Kernel80_Valid_Out, channel2_Kernel80_Valid_Out, channel3_Kernel80_Valid_Out, channel4_Kernel80_Valid_Out, channel5_Kernel80_Valid_Out, channel6_Kernel80_Valid_Out, channel7_Kernel80_Valid_Out, channel8_Kernel80_Valid_Out, channel9_Kernel80_Valid_Out, channel10_Kernel80_Valid_Out, channel11_Kernel80_Valid_Out, channel12_Kernel80_Valid_Out, channel13_Kernel80_Valid_Out, channel14_Kernel80_Valid_Out, channel15_Kernel80_Valid_Out, channel16_Kernel80_Valid_Out, channel17_Kernel80_Valid_Out, channel18_Kernel80_Valid_Out, channel19_Kernel80_Valid_Out, channel20_Kernel80_Valid_Out, channel21_Kernel80_Valid_Out, channel22_Kernel80_Valid_Out, channel23_Kernel80_Valid_Out, channel24_Kernel80_Valid_Out, channel25_Kernel80_Valid_Out, channel26_Kernel80_Valid_Out, channel27_Kernel80_Valid_Out, channel28_Kernel80_Valid_Out, channel29_Kernel80_Valid_Out, channel30_Kernel80_Valid_Out, channel31_Kernel80_Valid_Out, channel32_Kernel80_Valid_Out, channel33_Kernel80_Valid_Out, channel34_Kernel80_Valid_Out, channel35_Kernel80_Valid_Out, channel36_Kernel80_Valid_Out, channel37_Kernel80_Valid_Out, channel38_Kernel80_Valid_Out, channel39_Kernel80_Valid_Out, channel40_Kernel80_Valid_Out, channel41_Kernel80_Valid_Out, channel42_Kernel80_Valid_Out, channel43_Kernel80_Valid_Out, channel44_Kernel80_Valid_Out, channel45_Kernel80_Valid_Out, channel46_Kernel80_Valid_Out, channel47_Kernel80_Valid_Out, channel48_Kernel80_Valid_Out, channel49_Kernel80_Valid_Out, channel50_Kernel80_Valid_Out, channel51_Kernel80_Valid_Out, channel52_Kernel80_Valid_Out, channel53_Kernel80_Valid_Out, channel54_Kernel80_Valid_Out, channel55_Kernel80_Valid_Out, channel56_Kernel80_Valid_Out, channel57_Kernel80_Valid_Out, channel58_Kernel80_Valid_Out, channel59_Kernel80_Valid_Out, channel60_Kernel80_Valid_Out, channel61_Kernel80_Valid_Out, channel62_Kernel80_Valid_Out, channel63_Kernel80_Valid_Out, channel64_Kernel80_Valid_Out;

	assign add_kernel80=channel1_Kernel80_Valid_Out & channel2_Kernel80_Valid_Out & channel3_Kernel80_Valid_Out & channel4_Kernel80_Valid_Out & channel5_Kernel80_Valid_Out & channel6_Kernel80_Valid_Out & channel7_Kernel80_Valid_Out & channel8_Kernel80_Valid_Out & channel9_Kernel80_Valid_Out & channel10_Kernel80_Valid_Out & channel11_Kernel80_Valid_Out & channel12_Kernel80_Valid_Out & channel13_Kernel80_Valid_Out & channel14_Kernel80_Valid_Out & channel15_Kernel80_Valid_Out & channel16_Kernel80_Valid_Out & channel17_Kernel80_Valid_Out & channel18_Kernel80_Valid_Out & channel19_Kernel80_Valid_Out & channel20_Kernel80_Valid_Out & channel21_Kernel80_Valid_Out & channel22_Kernel80_Valid_Out & channel23_Kernel80_Valid_Out & channel24_Kernel80_Valid_Out & channel25_Kernel80_Valid_Out & channel26_Kernel80_Valid_Out & channel27_Kernel80_Valid_Out & channel28_Kernel80_Valid_Out & channel29_Kernel80_Valid_Out & channel30_Kernel80_Valid_Out & channel31_Kernel80_Valid_Out & channel32_Kernel80_Valid_Out & channel33_Kernel80_Valid_Out & channel34_Kernel80_Valid_Out & channel35_Kernel80_Valid_Out & channel36_Kernel80_Valid_Out & channel37_Kernel80_Valid_Out & channel38_Kernel80_Valid_Out & channel39_Kernel80_Valid_Out & channel40_Kernel80_Valid_Out & channel41_Kernel80_Valid_Out & channel42_Kernel80_Valid_Out & channel43_Kernel80_Valid_Out & channel44_Kernel80_Valid_Out & channel45_Kernel80_Valid_Out & channel46_Kernel80_Valid_Out & channel47_Kernel80_Valid_Out & channel48_Kernel80_Valid_Out & channel49_Kernel80_Valid_Out & channel50_Kernel80_Valid_Out & channel51_Kernel80_Valid_Out & channel52_Kernel80_Valid_Out & channel53_Kernel80_Valid_Out & channel54_Kernel80_Valid_Out & channel55_Kernel80_Valid_Out & channel56_Kernel80_Valid_Out & channel57_Kernel80_Valid_Out & channel58_Kernel80_Valid_Out & channel59_Kernel80_Valid_Out & channel60_Kernel80_Valid_Out & channel61_Kernel80_Valid_Out & channel62_Kernel80_Valid_Out & channel63_Kernel80_Valid_Out & channel64_Kernel80_Valid_Out;

	wire channel1_Kernel81_Valid_Out, channel2_Kernel81_Valid_Out, channel3_Kernel81_Valid_Out, channel4_Kernel81_Valid_Out, channel5_Kernel81_Valid_Out, channel6_Kernel81_Valid_Out, channel7_Kernel81_Valid_Out, channel8_Kernel81_Valid_Out, channel9_Kernel81_Valid_Out, channel10_Kernel81_Valid_Out, channel11_Kernel81_Valid_Out, channel12_Kernel81_Valid_Out, channel13_Kernel81_Valid_Out, channel14_Kernel81_Valid_Out, channel15_Kernel81_Valid_Out, channel16_Kernel81_Valid_Out, channel17_Kernel81_Valid_Out, channel18_Kernel81_Valid_Out, channel19_Kernel81_Valid_Out, channel20_Kernel81_Valid_Out, channel21_Kernel81_Valid_Out, channel22_Kernel81_Valid_Out, channel23_Kernel81_Valid_Out, channel24_Kernel81_Valid_Out, channel25_Kernel81_Valid_Out, channel26_Kernel81_Valid_Out, channel27_Kernel81_Valid_Out, channel28_Kernel81_Valid_Out, channel29_Kernel81_Valid_Out, channel30_Kernel81_Valid_Out, channel31_Kernel81_Valid_Out, channel32_Kernel81_Valid_Out, channel33_Kernel81_Valid_Out, channel34_Kernel81_Valid_Out, channel35_Kernel81_Valid_Out, channel36_Kernel81_Valid_Out, channel37_Kernel81_Valid_Out, channel38_Kernel81_Valid_Out, channel39_Kernel81_Valid_Out, channel40_Kernel81_Valid_Out, channel41_Kernel81_Valid_Out, channel42_Kernel81_Valid_Out, channel43_Kernel81_Valid_Out, channel44_Kernel81_Valid_Out, channel45_Kernel81_Valid_Out, channel46_Kernel81_Valid_Out, channel47_Kernel81_Valid_Out, channel48_Kernel81_Valid_Out, channel49_Kernel81_Valid_Out, channel50_Kernel81_Valid_Out, channel51_Kernel81_Valid_Out, channel52_Kernel81_Valid_Out, channel53_Kernel81_Valid_Out, channel54_Kernel81_Valid_Out, channel55_Kernel81_Valid_Out, channel56_Kernel81_Valid_Out, channel57_Kernel81_Valid_Out, channel58_Kernel81_Valid_Out, channel59_Kernel81_Valid_Out, channel60_Kernel81_Valid_Out, channel61_Kernel81_Valid_Out, channel62_Kernel81_Valid_Out, channel63_Kernel81_Valid_Out, channel64_Kernel81_Valid_Out;

	assign add_kernel81=channel1_Kernel81_Valid_Out & channel2_Kernel81_Valid_Out & channel3_Kernel81_Valid_Out & channel4_Kernel81_Valid_Out & channel5_Kernel81_Valid_Out & channel6_Kernel81_Valid_Out & channel7_Kernel81_Valid_Out & channel8_Kernel81_Valid_Out & channel9_Kernel81_Valid_Out & channel10_Kernel81_Valid_Out & channel11_Kernel81_Valid_Out & channel12_Kernel81_Valid_Out & channel13_Kernel81_Valid_Out & channel14_Kernel81_Valid_Out & channel15_Kernel81_Valid_Out & channel16_Kernel81_Valid_Out & channel17_Kernel81_Valid_Out & channel18_Kernel81_Valid_Out & channel19_Kernel81_Valid_Out & channel20_Kernel81_Valid_Out & channel21_Kernel81_Valid_Out & channel22_Kernel81_Valid_Out & channel23_Kernel81_Valid_Out & channel24_Kernel81_Valid_Out & channel25_Kernel81_Valid_Out & channel26_Kernel81_Valid_Out & channel27_Kernel81_Valid_Out & channel28_Kernel81_Valid_Out & channel29_Kernel81_Valid_Out & channel30_Kernel81_Valid_Out & channel31_Kernel81_Valid_Out & channel32_Kernel81_Valid_Out & channel33_Kernel81_Valid_Out & channel34_Kernel81_Valid_Out & channel35_Kernel81_Valid_Out & channel36_Kernel81_Valid_Out & channel37_Kernel81_Valid_Out & channel38_Kernel81_Valid_Out & channel39_Kernel81_Valid_Out & channel40_Kernel81_Valid_Out & channel41_Kernel81_Valid_Out & channel42_Kernel81_Valid_Out & channel43_Kernel81_Valid_Out & channel44_Kernel81_Valid_Out & channel45_Kernel81_Valid_Out & channel46_Kernel81_Valid_Out & channel47_Kernel81_Valid_Out & channel48_Kernel81_Valid_Out & channel49_Kernel81_Valid_Out & channel50_Kernel81_Valid_Out & channel51_Kernel81_Valid_Out & channel52_Kernel81_Valid_Out & channel53_Kernel81_Valid_Out & channel54_Kernel81_Valid_Out & channel55_Kernel81_Valid_Out & channel56_Kernel81_Valid_Out & channel57_Kernel81_Valid_Out & channel58_Kernel81_Valid_Out & channel59_Kernel81_Valid_Out & channel60_Kernel81_Valid_Out & channel61_Kernel81_Valid_Out & channel62_Kernel81_Valid_Out & channel63_Kernel81_Valid_Out & channel64_Kernel81_Valid_Out;

	wire channel1_Kernel82_Valid_Out, channel2_Kernel82_Valid_Out, channel3_Kernel82_Valid_Out, channel4_Kernel82_Valid_Out, channel5_Kernel82_Valid_Out, channel6_Kernel82_Valid_Out, channel7_Kernel82_Valid_Out, channel8_Kernel82_Valid_Out, channel9_Kernel82_Valid_Out, channel10_Kernel82_Valid_Out, channel11_Kernel82_Valid_Out, channel12_Kernel82_Valid_Out, channel13_Kernel82_Valid_Out, channel14_Kernel82_Valid_Out, channel15_Kernel82_Valid_Out, channel16_Kernel82_Valid_Out, channel17_Kernel82_Valid_Out, channel18_Kernel82_Valid_Out, channel19_Kernel82_Valid_Out, channel20_Kernel82_Valid_Out, channel21_Kernel82_Valid_Out, channel22_Kernel82_Valid_Out, channel23_Kernel82_Valid_Out, channel24_Kernel82_Valid_Out, channel25_Kernel82_Valid_Out, channel26_Kernel82_Valid_Out, channel27_Kernel82_Valid_Out, channel28_Kernel82_Valid_Out, channel29_Kernel82_Valid_Out, channel30_Kernel82_Valid_Out, channel31_Kernel82_Valid_Out, channel32_Kernel82_Valid_Out, channel33_Kernel82_Valid_Out, channel34_Kernel82_Valid_Out, channel35_Kernel82_Valid_Out, channel36_Kernel82_Valid_Out, channel37_Kernel82_Valid_Out, channel38_Kernel82_Valid_Out, channel39_Kernel82_Valid_Out, channel40_Kernel82_Valid_Out, channel41_Kernel82_Valid_Out, channel42_Kernel82_Valid_Out, channel43_Kernel82_Valid_Out, channel44_Kernel82_Valid_Out, channel45_Kernel82_Valid_Out, channel46_Kernel82_Valid_Out, channel47_Kernel82_Valid_Out, channel48_Kernel82_Valid_Out, channel49_Kernel82_Valid_Out, channel50_Kernel82_Valid_Out, channel51_Kernel82_Valid_Out, channel52_Kernel82_Valid_Out, channel53_Kernel82_Valid_Out, channel54_Kernel82_Valid_Out, channel55_Kernel82_Valid_Out, channel56_Kernel82_Valid_Out, channel57_Kernel82_Valid_Out, channel58_Kernel82_Valid_Out, channel59_Kernel82_Valid_Out, channel60_Kernel82_Valid_Out, channel61_Kernel82_Valid_Out, channel62_Kernel82_Valid_Out, channel63_Kernel82_Valid_Out, channel64_Kernel82_Valid_Out;

	assign add_kernel82=channel1_Kernel82_Valid_Out & channel2_Kernel82_Valid_Out & channel3_Kernel82_Valid_Out & channel4_Kernel82_Valid_Out & channel5_Kernel82_Valid_Out & channel6_Kernel82_Valid_Out & channel7_Kernel82_Valid_Out & channel8_Kernel82_Valid_Out & channel9_Kernel82_Valid_Out & channel10_Kernel82_Valid_Out & channel11_Kernel82_Valid_Out & channel12_Kernel82_Valid_Out & channel13_Kernel82_Valid_Out & channel14_Kernel82_Valid_Out & channel15_Kernel82_Valid_Out & channel16_Kernel82_Valid_Out & channel17_Kernel82_Valid_Out & channel18_Kernel82_Valid_Out & channel19_Kernel82_Valid_Out & channel20_Kernel82_Valid_Out & channel21_Kernel82_Valid_Out & channel22_Kernel82_Valid_Out & channel23_Kernel82_Valid_Out & channel24_Kernel82_Valid_Out & channel25_Kernel82_Valid_Out & channel26_Kernel82_Valid_Out & channel27_Kernel82_Valid_Out & channel28_Kernel82_Valid_Out & channel29_Kernel82_Valid_Out & channel30_Kernel82_Valid_Out & channel31_Kernel82_Valid_Out & channel32_Kernel82_Valid_Out & channel33_Kernel82_Valid_Out & channel34_Kernel82_Valid_Out & channel35_Kernel82_Valid_Out & channel36_Kernel82_Valid_Out & channel37_Kernel82_Valid_Out & channel38_Kernel82_Valid_Out & channel39_Kernel82_Valid_Out & channel40_Kernel82_Valid_Out & channel41_Kernel82_Valid_Out & channel42_Kernel82_Valid_Out & channel43_Kernel82_Valid_Out & channel44_Kernel82_Valid_Out & channel45_Kernel82_Valid_Out & channel46_Kernel82_Valid_Out & channel47_Kernel82_Valid_Out & channel48_Kernel82_Valid_Out & channel49_Kernel82_Valid_Out & channel50_Kernel82_Valid_Out & channel51_Kernel82_Valid_Out & channel52_Kernel82_Valid_Out & channel53_Kernel82_Valid_Out & channel54_Kernel82_Valid_Out & channel55_Kernel82_Valid_Out & channel56_Kernel82_Valid_Out & channel57_Kernel82_Valid_Out & channel58_Kernel82_Valid_Out & channel59_Kernel82_Valid_Out & channel60_Kernel82_Valid_Out & channel61_Kernel82_Valid_Out & channel62_Kernel82_Valid_Out & channel63_Kernel82_Valid_Out & channel64_Kernel82_Valid_Out;

	wire channel1_Kernel83_Valid_Out, channel2_Kernel83_Valid_Out, channel3_Kernel83_Valid_Out, channel4_Kernel83_Valid_Out, channel5_Kernel83_Valid_Out, channel6_Kernel83_Valid_Out, channel7_Kernel83_Valid_Out, channel8_Kernel83_Valid_Out, channel9_Kernel83_Valid_Out, channel10_Kernel83_Valid_Out, channel11_Kernel83_Valid_Out, channel12_Kernel83_Valid_Out, channel13_Kernel83_Valid_Out, channel14_Kernel83_Valid_Out, channel15_Kernel83_Valid_Out, channel16_Kernel83_Valid_Out, channel17_Kernel83_Valid_Out, channel18_Kernel83_Valid_Out, channel19_Kernel83_Valid_Out, channel20_Kernel83_Valid_Out, channel21_Kernel83_Valid_Out, channel22_Kernel83_Valid_Out, channel23_Kernel83_Valid_Out, channel24_Kernel83_Valid_Out, channel25_Kernel83_Valid_Out, channel26_Kernel83_Valid_Out, channel27_Kernel83_Valid_Out, channel28_Kernel83_Valid_Out, channel29_Kernel83_Valid_Out, channel30_Kernel83_Valid_Out, channel31_Kernel83_Valid_Out, channel32_Kernel83_Valid_Out, channel33_Kernel83_Valid_Out, channel34_Kernel83_Valid_Out, channel35_Kernel83_Valid_Out, channel36_Kernel83_Valid_Out, channel37_Kernel83_Valid_Out, channel38_Kernel83_Valid_Out, channel39_Kernel83_Valid_Out, channel40_Kernel83_Valid_Out, channel41_Kernel83_Valid_Out, channel42_Kernel83_Valid_Out, channel43_Kernel83_Valid_Out, channel44_Kernel83_Valid_Out, channel45_Kernel83_Valid_Out, channel46_Kernel83_Valid_Out, channel47_Kernel83_Valid_Out, channel48_Kernel83_Valid_Out, channel49_Kernel83_Valid_Out, channel50_Kernel83_Valid_Out, channel51_Kernel83_Valid_Out, channel52_Kernel83_Valid_Out, channel53_Kernel83_Valid_Out, channel54_Kernel83_Valid_Out, channel55_Kernel83_Valid_Out, channel56_Kernel83_Valid_Out, channel57_Kernel83_Valid_Out, channel58_Kernel83_Valid_Out, channel59_Kernel83_Valid_Out, channel60_Kernel83_Valid_Out, channel61_Kernel83_Valid_Out, channel62_Kernel83_Valid_Out, channel63_Kernel83_Valid_Out, channel64_Kernel83_Valid_Out;

	assign add_kernel83=channel1_Kernel83_Valid_Out & channel2_Kernel83_Valid_Out & channel3_Kernel83_Valid_Out & channel4_Kernel83_Valid_Out & channel5_Kernel83_Valid_Out & channel6_Kernel83_Valid_Out & channel7_Kernel83_Valid_Out & channel8_Kernel83_Valid_Out & channel9_Kernel83_Valid_Out & channel10_Kernel83_Valid_Out & channel11_Kernel83_Valid_Out & channel12_Kernel83_Valid_Out & channel13_Kernel83_Valid_Out & channel14_Kernel83_Valid_Out & channel15_Kernel83_Valid_Out & channel16_Kernel83_Valid_Out & channel17_Kernel83_Valid_Out & channel18_Kernel83_Valid_Out & channel19_Kernel83_Valid_Out & channel20_Kernel83_Valid_Out & channel21_Kernel83_Valid_Out & channel22_Kernel83_Valid_Out & channel23_Kernel83_Valid_Out & channel24_Kernel83_Valid_Out & channel25_Kernel83_Valid_Out & channel26_Kernel83_Valid_Out & channel27_Kernel83_Valid_Out & channel28_Kernel83_Valid_Out & channel29_Kernel83_Valid_Out & channel30_Kernel83_Valid_Out & channel31_Kernel83_Valid_Out & channel32_Kernel83_Valid_Out & channel33_Kernel83_Valid_Out & channel34_Kernel83_Valid_Out & channel35_Kernel83_Valid_Out & channel36_Kernel83_Valid_Out & channel37_Kernel83_Valid_Out & channel38_Kernel83_Valid_Out & channel39_Kernel83_Valid_Out & channel40_Kernel83_Valid_Out & channel41_Kernel83_Valid_Out & channel42_Kernel83_Valid_Out & channel43_Kernel83_Valid_Out & channel44_Kernel83_Valid_Out & channel45_Kernel83_Valid_Out & channel46_Kernel83_Valid_Out & channel47_Kernel83_Valid_Out & channel48_Kernel83_Valid_Out & channel49_Kernel83_Valid_Out & channel50_Kernel83_Valid_Out & channel51_Kernel83_Valid_Out & channel52_Kernel83_Valid_Out & channel53_Kernel83_Valid_Out & channel54_Kernel83_Valid_Out & channel55_Kernel83_Valid_Out & channel56_Kernel83_Valid_Out & channel57_Kernel83_Valid_Out & channel58_Kernel83_Valid_Out & channel59_Kernel83_Valid_Out & channel60_Kernel83_Valid_Out & channel61_Kernel83_Valid_Out & channel62_Kernel83_Valid_Out & channel63_Kernel83_Valid_Out & channel64_Kernel83_Valid_Out;

	wire channel1_Kernel84_Valid_Out, channel2_Kernel84_Valid_Out, channel3_Kernel84_Valid_Out, channel4_Kernel84_Valid_Out, channel5_Kernel84_Valid_Out, channel6_Kernel84_Valid_Out, channel7_Kernel84_Valid_Out, channel8_Kernel84_Valid_Out, channel9_Kernel84_Valid_Out, channel10_Kernel84_Valid_Out, channel11_Kernel84_Valid_Out, channel12_Kernel84_Valid_Out, channel13_Kernel84_Valid_Out, channel14_Kernel84_Valid_Out, channel15_Kernel84_Valid_Out, channel16_Kernel84_Valid_Out, channel17_Kernel84_Valid_Out, channel18_Kernel84_Valid_Out, channel19_Kernel84_Valid_Out, channel20_Kernel84_Valid_Out, channel21_Kernel84_Valid_Out, channel22_Kernel84_Valid_Out, channel23_Kernel84_Valid_Out, channel24_Kernel84_Valid_Out, channel25_Kernel84_Valid_Out, channel26_Kernel84_Valid_Out, channel27_Kernel84_Valid_Out, channel28_Kernel84_Valid_Out, channel29_Kernel84_Valid_Out, channel30_Kernel84_Valid_Out, channel31_Kernel84_Valid_Out, channel32_Kernel84_Valid_Out, channel33_Kernel84_Valid_Out, channel34_Kernel84_Valid_Out, channel35_Kernel84_Valid_Out, channel36_Kernel84_Valid_Out, channel37_Kernel84_Valid_Out, channel38_Kernel84_Valid_Out, channel39_Kernel84_Valid_Out, channel40_Kernel84_Valid_Out, channel41_Kernel84_Valid_Out, channel42_Kernel84_Valid_Out, channel43_Kernel84_Valid_Out, channel44_Kernel84_Valid_Out, channel45_Kernel84_Valid_Out, channel46_Kernel84_Valid_Out, channel47_Kernel84_Valid_Out, channel48_Kernel84_Valid_Out, channel49_Kernel84_Valid_Out, channel50_Kernel84_Valid_Out, channel51_Kernel84_Valid_Out, channel52_Kernel84_Valid_Out, channel53_Kernel84_Valid_Out, channel54_Kernel84_Valid_Out, channel55_Kernel84_Valid_Out, channel56_Kernel84_Valid_Out, channel57_Kernel84_Valid_Out, channel58_Kernel84_Valid_Out, channel59_Kernel84_Valid_Out, channel60_Kernel84_Valid_Out, channel61_Kernel84_Valid_Out, channel62_Kernel84_Valid_Out, channel63_Kernel84_Valid_Out, channel64_Kernel84_Valid_Out;

	assign add_kernel84=channel1_Kernel84_Valid_Out & channel2_Kernel84_Valid_Out & channel3_Kernel84_Valid_Out & channel4_Kernel84_Valid_Out & channel5_Kernel84_Valid_Out & channel6_Kernel84_Valid_Out & channel7_Kernel84_Valid_Out & channel8_Kernel84_Valid_Out & channel9_Kernel84_Valid_Out & channel10_Kernel84_Valid_Out & channel11_Kernel84_Valid_Out & channel12_Kernel84_Valid_Out & channel13_Kernel84_Valid_Out & channel14_Kernel84_Valid_Out & channel15_Kernel84_Valid_Out & channel16_Kernel84_Valid_Out & channel17_Kernel84_Valid_Out & channel18_Kernel84_Valid_Out & channel19_Kernel84_Valid_Out & channel20_Kernel84_Valid_Out & channel21_Kernel84_Valid_Out & channel22_Kernel84_Valid_Out & channel23_Kernel84_Valid_Out & channel24_Kernel84_Valid_Out & channel25_Kernel84_Valid_Out & channel26_Kernel84_Valid_Out & channel27_Kernel84_Valid_Out & channel28_Kernel84_Valid_Out & channel29_Kernel84_Valid_Out & channel30_Kernel84_Valid_Out & channel31_Kernel84_Valid_Out & channel32_Kernel84_Valid_Out & channel33_Kernel84_Valid_Out & channel34_Kernel84_Valid_Out & channel35_Kernel84_Valid_Out & channel36_Kernel84_Valid_Out & channel37_Kernel84_Valid_Out & channel38_Kernel84_Valid_Out & channel39_Kernel84_Valid_Out & channel40_Kernel84_Valid_Out & channel41_Kernel84_Valid_Out & channel42_Kernel84_Valid_Out & channel43_Kernel84_Valid_Out & channel44_Kernel84_Valid_Out & channel45_Kernel84_Valid_Out & channel46_Kernel84_Valid_Out & channel47_Kernel84_Valid_Out & channel48_Kernel84_Valid_Out & channel49_Kernel84_Valid_Out & channel50_Kernel84_Valid_Out & channel51_Kernel84_Valid_Out & channel52_Kernel84_Valid_Out & channel53_Kernel84_Valid_Out & channel54_Kernel84_Valid_Out & channel55_Kernel84_Valid_Out & channel56_Kernel84_Valid_Out & channel57_Kernel84_Valid_Out & channel58_Kernel84_Valid_Out & channel59_Kernel84_Valid_Out & channel60_Kernel84_Valid_Out & channel61_Kernel84_Valid_Out & channel62_Kernel84_Valid_Out & channel63_Kernel84_Valid_Out & channel64_Kernel84_Valid_Out;

	wire channel1_Kernel85_Valid_Out, channel2_Kernel85_Valid_Out, channel3_Kernel85_Valid_Out, channel4_Kernel85_Valid_Out, channel5_Kernel85_Valid_Out, channel6_Kernel85_Valid_Out, channel7_Kernel85_Valid_Out, channel8_Kernel85_Valid_Out, channel9_Kernel85_Valid_Out, channel10_Kernel85_Valid_Out, channel11_Kernel85_Valid_Out, channel12_Kernel85_Valid_Out, channel13_Kernel85_Valid_Out, channel14_Kernel85_Valid_Out, channel15_Kernel85_Valid_Out, channel16_Kernel85_Valid_Out, channel17_Kernel85_Valid_Out, channel18_Kernel85_Valid_Out, channel19_Kernel85_Valid_Out, channel20_Kernel85_Valid_Out, channel21_Kernel85_Valid_Out, channel22_Kernel85_Valid_Out, channel23_Kernel85_Valid_Out, channel24_Kernel85_Valid_Out, channel25_Kernel85_Valid_Out, channel26_Kernel85_Valid_Out, channel27_Kernel85_Valid_Out, channel28_Kernel85_Valid_Out, channel29_Kernel85_Valid_Out, channel30_Kernel85_Valid_Out, channel31_Kernel85_Valid_Out, channel32_Kernel85_Valid_Out, channel33_Kernel85_Valid_Out, channel34_Kernel85_Valid_Out, channel35_Kernel85_Valid_Out, channel36_Kernel85_Valid_Out, channel37_Kernel85_Valid_Out, channel38_Kernel85_Valid_Out, channel39_Kernel85_Valid_Out, channel40_Kernel85_Valid_Out, channel41_Kernel85_Valid_Out, channel42_Kernel85_Valid_Out, channel43_Kernel85_Valid_Out, channel44_Kernel85_Valid_Out, channel45_Kernel85_Valid_Out, channel46_Kernel85_Valid_Out, channel47_Kernel85_Valid_Out, channel48_Kernel85_Valid_Out, channel49_Kernel85_Valid_Out, channel50_Kernel85_Valid_Out, channel51_Kernel85_Valid_Out, channel52_Kernel85_Valid_Out, channel53_Kernel85_Valid_Out, channel54_Kernel85_Valid_Out, channel55_Kernel85_Valid_Out, channel56_Kernel85_Valid_Out, channel57_Kernel85_Valid_Out, channel58_Kernel85_Valid_Out, channel59_Kernel85_Valid_Out, channel60_Kernel85_Valid_Out, channel61_Kernel85_Valid_Out, channel62_Kernel85_Valid_Out, channel63_Kernel85_Valid_Out, channel64_Kernel85_Valid_Out;

	assign add_kernel85=channel1_Kernel85_Valid_Out & channel2_Kernel85_Valid_Out & channel3_Kernel85_Valid_Out & channel4_Kernel85_Valid_Out & channel5_Kernel85_Valid_Out & channel6_Kernel85_Valid_Out & channel7_Kernel85_Valid_Out & channel8_Kernel85_Valid_Out & channel9_Kernel85_Valid_Out & channel10_Kernel85_Valid_Out & channel11_Kernel85_Valid_Out & channel12_Kernel85_Valid_Out & channel13_Kernel85_Valid_Out & channel14_Kernel85_Valid_Out & channel15_Kernel85_Valid_Out & channel16_Kernel85_Valid_Out & channel17_Kernel85_Valid_Out & channel18_Kernel85_Valid_Out & channel19_Kernel85_Valid_Out & channel20_Kernel85_Valid_Out & channel21_Kernel85_Valid_Out & channel22_Kernel85_Valid_Out & channel23_Kernel85_Valid_Out & channel24_Kernel85_Valid_Out & channel25_Kernel85_Valid_Out & channel26_Kernel85_Valid_Out & channel27_Kernel85_Valid_Out & channel28_Kernel85_Valid_Out & channel29_Kernel85_Valid_Out & channel30_Kernel85_Valid_Out & channel31_Kernel85_Valid_Out & channel32_Kernel85_Valid_Out & channel33_Kernel85_Valid_Out & channel34_Kernel85_Valid_Out & channel35_Kernel85_Valid_Out & channel36_Kernel85_Valid_Out & channel37_Kernel85_Valid_Out & channel38_Kernel85_Valid_Out & channel39_Kernel85_Valid_Out & channel40_Kernel85_Valid_Out & channel41_Kernel85_Valid_Out & channel42_Kernel85_Valid_Out & channel43_Kernel85_Valid_Out & channel44_Kernel85_Valid_Out & channel45_Kernel85_Valid_Out & channel46_Kernel85_Valid_Out & channel47_Kernel85_Valid_Out & channel48_Kernel85_Valid_Out & channel49_Kernel85_Valid_Out & channel50_Kernel85_Valid_Out & channel51_Kernel85_Valid_Out & channel52_Kernel85_Valid_Out & channel53_Kernel85_Valid_Out & channel54_Kernel85_Valid_Out & channel55_Kernel85_Valid_Out & channel56_Kernel85_Valid_Out & channel57_Kernel85_Valid_Out & channel58_Kernel85_Valid_Out & channel59_Kernel85_Valid_Out & channel60_Kernel85_Valid_Out & channel61_Kernel85_Valid_Out & channel62_Kernel85_Valid_Out & channel63_Kernel85_Valid_Out & channel64_Kernel85_Valid_Out;

	wire channel1_Kernel86_Valid_Out, channel2_Kernel86_Valid_Out, channel3_Kernel86_Valid_Out, channel4_Kernel86_Valid_Out, channel5_Kernel86_Valid_Out, channel6_Kernel86_Valid_Out, channel7_Kernel86_Valid_Out, channel8_Kernel86_Valid_Out, channel9_Kernel86_Valid_Out, channel10_Kernel86_Valid_Out, channel11_Kernel86_Valid_Out, channel12_Kernel86_Valid_Out, channel13_Kernel86_Valid_Out, channel14_Kernel86_Valid_Out, channel15_Kernel86_Valid_Out, channel16_Kernel86_Valid_Out, channel17_Kernel86_Valid_Out, channel18_Kernel86_Valid_Out, channel19_Kernel86_Valid_Out, channel20_Kernel86_Valid_Out, channel21_Kernel86_Valid_Out, channel22_Kernel86_Valid_Out, channel23_Kernel86_Valid_Out, channel24_Kernel86_Valid_Out, channel25_Kernel86_Valid_Out, channel26_Kernel86_Valid_Out, channel27_Kernel86_Valid_Out, channel28_Kernel86_Valid_Out, channel29_Kernel86_Valid_Out, channel30_Kernel86_Valid_Out, channel31_Kernel86_Valid_Out, channel32_Kernel86_Valid_Out, channel33_Kernel86_Valid_Out, channel34_Kernel86_Valid_Out, channel35_Kernel86_Valid_Out, channel36_Kernel86_Valid_Out, channel37_Kernel86_Valid_Out, channel38_Kernel86_Valid_Out, channel39_Kernel86_Valid_Out, channel40_Kernel86_Valid_Out, channel41_Kernel86_Valid_Out, channel42_Kernel86_Valid_Out, channel43_Kernel86_Valid_Out, channel44_Kernel86_Valid_Out, channel45_Kernel86_Valid_Out, channel46_Kernel86_Valid_Out, channel47_Kernel86_Valid_Out, channel48_Kernel86_Valid_Out, channel49_Kernel86_Valid_Out, channel50_Kernel86_Valid_Out, channel51_Kernel86_Valid_Out, channel52_Kernel86_Valid_Out, channel53_Kernel86_Valid_Out, channel54_Kernel86_Valid_Out, channel55_Kernel86_Valid_Out, channel56_Kernel86_Valid_Out, channel57_Kernel86_Valid_Out, channel58_Kernel86_Valid_Out, channel59_Kernel86_Valid_Out, channel60_Kernel86_Valid_Out, channel61_Kernel86_Valid_Out, channel62_Kernel86_Valid_Out, channel63_Kernel86_Valid_Out, channel64_Kernel86_Valid_Out;

	assign add_kernel86=channel1_Kernel86_Valid_Out & channel2_Kernel86_Valid_Out & channel3_Kernel86_Valid_Out & channel4_Kernel86_Valid_Out & channel5_Kernel86_Valid_Out & channel6_Kernel86_Valid_Out & channel7_Kernel86_Valid_Out & channel8_Kernel86_Valid_Out & channel9_Kernel86_Valid_Out & channel10_Kernel86_Valid_Out & channel11_Kernel86_Valid_Out & channel12_Kernel86_Valid_Out & channel13_Kernel86_Valid_Out & channel14_Kernel86_Valid_Out & channel15_Kernel86_Valid_Out & channel16_Kernel86_Valid_Out & channel17_Kernel86_Valid_Out & channel18_Kernel86_Valid_Out & channel19_Kernel86_Valid_Out & channel20_Kernel86_Valid_Out & channel21_Kernel86_Valid_Out & channel22_Kernel86_Valid_Out & channel23_Kernel86_Valid_Out & channel24_Kernel86_Valid_Out & channel25_Kernel86_Valid_Out & channel26_Kernel86_Valid_Out & channel27_Kernel86_Valid_Out & channel28_Kernel86_Valid_Out & channel29_Kernel86_Valid_Out & channel30_Kernel86_Valid_Out & channel31_Kernel86_Valid_Out & channel32_Kernel86_Valid_Out & channel33_Kernel86_Valid_Out & channel34_Kernel86_Valid_Out & channel35_Kernel86_Valid_Out & channel36_Kernel86_Valid_Out & channel37_Kernel86_Valid_Out & channel38_Kernel86_Valid_Out & channel39_Kernel86_Valid_Out & channel40_Kernel86_Valid_Out & channel41_Kernel86_Valid_Out & channel42_Kernel86_Valid_Out & channel43_Kernel86_Valid_Out & channel44_Kernel86_Valid_Out & channel45_Kernel86_Valid_Out & channel46_Kernel86_Valid_Out & channel47_Kernel86_Valid_Out & channel48_Kernel86_Valid_Out & channel49_Kernel86_Valid_Out & channel50_Kernel86_Valid_Out & channel51_Kernel86_Valid_Out & channel52_Kernel86_Valid_Out & channel53_Kernel86_Valid_Out & channel54_Kernel86_Valid_Out & channel55_Kernel86_Valid_Out & channel56_Kernel86_Valid_Out & channel57_Kernel86_Valid_Out & channel58_Kernel86_Valid_Out & channel59_Kernel86_Valid_Out & channel60_Kernel86_Valid_Out & channel61_Kernel86_Valid_Out & channel62_Kernel86_Valid_Out & channel63_Kernel86_Valid_Out & channel64_Kernel86_Valid_Out;

	wire channel1_Kernel87_Valid_Out, channel2_Kernel87_Valid_Out, channel3_Kernel87_Valid_Out, channel4_Kernel87_Valid_Out, channel5_Kernel87_Valid_Out, channel6_Kernel87_Valid_Out, channel7_Kernel87_Valid_Out, channel8_Kernel87_Valid_Out, channel9_Kernel87_Valid_Out, channel10_Kernel87_Valid_Out, channel11_Kernel87_Valid_Out, channel12_Kernel87_Valid_Out, channel13_Kernel87_Valid_Out, channel14_Kernel87_Valid_Out, channel15_Kernel87_Valid_Out, channel16_Kernel87_Valid_Out, channel17_Kernel87_Valid_Out, channel18_Kernel87_Valid_Out, channel19_Kernel87_Valid_Out, channel20_Kernel87_Valid_Out, channel21_Kernel87_Valid_Out, channel22_Kernel87_Valid_Out, channel23_Kernel87_Valid_Out, channel24_Kernel87_Valid_Out, channel25_Kernel87_Valid_Out, channel26_Kernel87_Valid_Out, channel27_Kernel87_Valid_Out, channel28_Kernel87_Valid_Out, channel29_Kernel87_Valid_Out, channel30_Kernel87_Valid_Out, channel31_Kernel87_Valid_Out, channel32_Kernel87_Valid_Out, channel33_Kernel87_Valid_Out, channel34_Kernel87_Valid_Out, channel35_Kernel87_Valid_Out, channel36_Kernel87_Valid_Out, channel37_Kernel87_Valid_Out, channel38_Kernel87_Valid_Out, channel39_Kernel87_Valid_Out, channel40_Kernel87_Valid_Out, channel41_Kernel87_Valid_Out, channel42_Kernel87_Valid_Out, channel43_Kernel87_Valid_Out, channel44_Kernel87_Valid_Out, channel45_Kernel87_Valid_Out, channel46_Kernel87_Valid_Out, channel47_Kernel87_Valid_Out, channel48_Kernel87_Valid_Out, channel49_Kernel87_Valid_Out, channel50_Kernel87_Valid_Out, channel51_Kernel87_Valid_Out, channel52_Kernel87_Valid_Out, channel53_Kernel87_Valid_Out, channel54_Kernel87_Valid_Out, channel55_Kernel87_Valid_Out, channel56_Kernel87_Valid_Out, channel57_Kernel87_Valid_Out, channel58_Kernel87_Valid_Out, channel59_Kernel87_Valid_Out, channel60_Kernel87_Valid_Out, channel61_Kernel87_Valid_Out, channel62_Kernel87_Valid_Out, channel63_Kernel87_Valid_Out, channel64_Kernel87_Valid_Out;

	assign add_kernel87=channel1_Kernel87_Valid_Out & channel2_Kernel87_Valid_Out & channel3_Kernel87_Valid_Out & channel4_Kernel87_Valid_Out & channel5_Kernel87_Valid_Out & channel6_Kernel87_Valid_Out & channel7_Kernel87_Valid_Out & channel8_Kernel87_Valid_Out & channel9_Kernel87_Valid_Out & channel10_Kernel87_Valid_Out & channel11_Kernel87_Valid_Out & channel12_Kernel87_Valid_Out & channel13_Kernel87_Valid_Out & channel14_Kernel87_Valid_Out & channel15_Kernel87_Valid_Out & channel16_Kernel87_Valid_Out & channel17_Kernel87_Valid_Out & channel18_Kernel87_Valid_Out & channel19_Kernel87_Valid_Out & channel20_Kernel87_Valid_Out & channel21_Kernel87_Valid_Out & channel22_Kernel87_Valid_Out & channel23_Kernel87_Valid_Out & channel24_Kernel87_Valid_Out & channel25_Kernel87_Valid_Out & channel26_Kernel87_Valid_Out & channel27_Kernel87_Valid_Out & channel28_Kernel87_Valid_Out & channel29_Kernel87_Valid_Out & channel30_Kernel87_Valid_Out & channel31_Kernel87_Valid_Out & channel32_Kernel87_Valid_Out & channel33_Kernel87_Valid_Out & channel34_Kernel87_Valid_Out & channel35_Kernel87_Valid_Out & channel36_Kernel87_Valid_Out & channel37_Kernel87_Valid_Out & channel38_Kernel87_Valid_Out & channel39_Kernel87_Valid_Out & channel40_Kernel87_Valid_Out & channel41_Kernel87_Valid_Out & channel42_Kernel87_Valid_Out & channel43_Kernel87_Valid_Out & channel44_Kernel87_Valid_Out & channel45_Kernel87_Valid_Out & channel46_Kernel87_Valid_Out & channel47_Kernel87_Valid_Out & channel48_Kernel87_Valid_Out & channel49_Kernel87_Valid_Out & channel50_Kernel87_Valid_Out & channel51_Kernel87_Valid_Out & channel52_Kernel87_Valid_Out & channel53_Kernel87_Valid_Out & channel54_Kernel87_Valid_Out & channel55_Kernel87_Valid_Out & channel56_Kernel87_Valid_Out & channel57_Kernel87_Valid_Out & channel58_Kernel87_Valid_Out & channel59_Kernel87_Valid_Out & channel60_Kernel87_Valid_Out & channel61_Kernel87_Valid_Out & channel62_Kernel87_Valid_Out & channel63_Kernel87_Valid_Out & channel64_Kernel87_Valid_Out;

	wire channel1_Kernel88_Valid_Out, channel2_Kernel88_Valid_Out, channel3_Kernel88_Valid_Out, channel4_Kernel88_Valid_Out, channel5_Kernel88_Valid_Out, channel6_Kernel88_Valid_Out, channel7_Kernel88_Valid_Out, channel8_Kernel88_Valid_Out, channel9_Kernel88_Valid_Out, channel10_Kernel88_Valid_Out, channel11_Kernel88_Valid_Out, channel12_Kernel88_Valid_Out, channel13_Kernel88_Valid_Out, channel14_Kernel88_Valid_Out, channel15_Kernel88_Valid_Out, channel16_Kernel88_Valid_Out, channel17_Kernel88_Valid_Out, channel18_Kernel88_Valid_Out, channel19_Kernel88_Valid_Out, channel20_Kernel88_Valid_Out, channel21_Kernel88_Valid_Out, channel22_Kernel88_Valid_Out, channel23_Kernel88_Valid_Out, channel24_Kernel88_Valid_Out, channel25_Kernel88_Valid_Out, channel26_Kernel88_Valid_Out, channel27_Kernel88_Valid_Out, channel28_Kernel88_Valid_Out, channel29_Kernel88_Valid_Out, channel30_Kernel88_Valid_Out, channel31_Kernel88_Valid_Out, channel32_Kernel88_Valid_Out, channel33_Kernel88_Valid_Out, channel34_Kernel88_Valid_Out, channel35_Kernel88_Valid_Out, channel36_Kernel88_Valid_Out, channel37_Kernel88_Valid_Out, channel38_Kernel88_Valid_Out, channel39_Kernel88_Valid_Out, channel40_Kernel88_Valid_Out, channel41_Kernel88_Valid_Out, channel42_Kernel88_Valid_Out, channel43_Kernel88_Valid_Out, channel44_Kernel88_Valid_Out, channel45_Kernel88_Valid_Out, channel46_Kernel88_Valid_Out, channel47_Kernel88_Valid_Out, channel48_Kernel88_Valid_Out, channel49_Kernel88_Valid_Out, channel50_Kernel88_Valid_Out, channel51_Kernel88_Valid_Out, channel52_Kernel88_Valid_Out, channel53_Kernel88_Valid_Out, channel54_Kernel88_Valid_Out, channel55_Kernel88_Valid_Out, channel56_Kernel88_Valid_Out, channel57_Kernel88_Valid_Out, channel58_Kernel88_Valid_Out, channel59_Kernel88_Valid_Out, channel60_Kernel88_Valid_Out, channel61_Kernel88_Valid_Out, channel62_Kernel88_Valid_Out, channel63_Kernel88_Valid_Out, channel64_Kernel88_Valid_Out;

	assign add_kernel88=channel1_Kernel88_Valid_Out & channel2_Kernel88_Valid_Out & channel3_Kernel88_Valid_Out & channel4_Kernel88_Valid_Out & channel5_Kernel88_Valid_Out & channel6_Kernel88_Valid_Out & channel7_Kernel88_Valid_Out & channel8_Kernel88_Valid_Out & channel9_Kernel88_Valid_Out & channel10_Kernel88_Valid_Out & channel11_Kernel88_Valid_Out & channel12_Kernel88_Valid_Out & channel13_Kernel88_Valid_Out & channel14_Kernel88_Valid_Out & channel15_Kernel88_Valid_Out & channel16_Kernel88_Valid_Out & channel17_Kernel88_Valid_Out & channel18_Kernel88_Valid_Out & channel19_Kernel88_Valid_Out & channel20_Kernel88_Valid_Out & channel21_Kernel88_Valid_Out & channel22_Kernel88_Valid_Out & channel23_Kernel88_Valid_Out & channel24_Kernel88_Valid_Out & channel25_Kernel88_Valid_Out & channel26_Kernel88_Valid_Out & channel27_Kernel88_Valid_Out & channel28_Kernel88_Valid_Out & channel29_Kernel88_Valid_Out & channel30_Kernel88_Valid_Out & channel31_Kernel88_Valid_Out & channel32_Kernel88_Valid_Out & channel33_Kernel88_Valid_Out & channel34_Kernel88_Valid_Out & channel35_Kernel88_Valid_Out & channel36_Kernel88_Valid_Out & channel37_Kernel88_Valid_Out & channel38_Kernel88_Valid_Out & channel39_Kernel88_Valid_Out & channel40_Kernel88_Valid_Out & channel41_Kernel88_Valid_Out & channel42_Kernel88_Valid_Out & channel43_Kernel88_Valid_Out & channel44_Kernel88_Valid_Out & channel45_Kernel88_Valid_Out & channel46_Kernel88_Valid_Out & channel47_Kernel88_Valid_Out & channel48_Kernel88_Valid_Out & channel49_Kernel88_Valid_Out & channel50_Kernel88_Valid_Out & channel51_Kernel88_Valid_Out & channel52_Kernel88_Valid_Out & channel53_Kernel88_Valid_Out & channel54_Kernel88_Valid_Out & channel55_Kernel88_Valid_Out & channel56_Kernel88_Valid_Out & channel57_Kernel88_Valid_Out & channel58_Kernel88_Valid_Out & channel59_Kernel88_Valid_Out & channel60_Kernel88_Valid_Out & channel61_Kernel88_Valid_Out & channel62_Kernel88_Valid_Out & channel63_Kernel88_Valid_Out & channel64_Kernel88_Valid_Out;

	wire channel1_Kernel89_Valid_Out, channel2_Kernel89_Valid_Out, channel3_Kernel89_Valid_Out, channel4_Kernel89_Valid_Out, channel5_Kernel89_Valid_Out, channel6_Kernel89_Valid_Out, channel7_Kernel89_Valid_Out, channel8_Kernel89_Valid_Out, channel9_Kernel89_Valid_Out, channel10_Kernel89_Valid_Out, channel11_Kernel89_Valid_Out, channel12_Kernel89_Valid_Out, channel13_Kernel89_Valid_Out, channel14_Kernel89_Valid_Out, channel15_Kernel89_Valid_Out, channel16_Kernel89_Valid_Out, channel17_Kernel89_Valid_Out, channel18_Kernel89_Valid_Out, channel19_Kernel89_Valid_Out, channel20_Kernel89_Valid_Out, channel21_Kernel89_Valid_Out, channel22_Kernel89_Valid_Out, channel23_Kernel89_Valid_Out, channel24_Kernel89_Valid_Out, channel25_Kernel89_Valid_Out, channel26_Kernel89_Valid_Out, channel27_Kernel89_Valid_Out, channel28_Kernel89_Valid_Out, channel29_Kernel89_Valid_Out, channel30_Kernel89_Valid_Out, channel31_Kernel89_Valid_Out, channel32_Kernel89_Valid_Out, channel33_Kernel89_Valid_Out, channel34_Kernel89_Valid_Out, channel35_Kernel89_Valid_Out, channel36_Kernel89_Valid_Out, channel37_Kernel89_Valid_Out, channel38_Kernel89_Valid_Out, channel39_Kernel89_Valid_Out, channel40_Kernel89_Valid_Out, channel41_Kernel89_Valid_Out, channel42_Kernel89_Valid_Out, channel43_Kernel89_Valid_Out, channel44_Kernel89_Valid_Out, channel45_Kernel89_Valid_Out, channel46_Kernel89_Valid_Out, channel47_Kernel89_Valid_Out, channel48_Kernel89_Valid_Out, channel49_Kernel89_Valid_Out, channel50_Kernel89_Valid_Out, channel51_Kernel89_Valid_Out, channel52_Kernel89_Valid_Out, channel53_Kernel89_Valid_Out, channel54_Kernel89_Valid_Out, channel55_Kernel89_Valid_Out, channel56_Kernel89_Valid_Out, channel57_Kernel89_Valid_Out, channel58_Kernel89_Valid_Out, channel59_Kernel89_Valid_Out, channel60_Kernel89_Valid_Out, channel61_Kernel89_Valid_Out, channel62_Kernel89_Valid_Out, channel63_Kernel89_Valid_Out, channel64_Kernel89_Valid_Out;

	assign add_kernel89=channel1_Kernel89_Valid_Out & channel2_Kernel89_Valid_Out & channel3_Kernel89_Valid_Out & channel4_Kernel89_Valid_Out & channel5_Kernel89_Valid_Out & channel6_Kernel89_Valid_Out & channel7_Kernel89_Valid_Out & channel8_Kernel89_Valid_Out & channel9_Kernel89_Valid_Out & channel10_Kernel89_Valid_Out & channel11_Kernel89_Valid_Out & channel12_Kernel89_Valid_Out & channel13_Kernel89_Valid_Out & channel14_Kernel89_Valid_Out & channel15_Kernel89_Valid_Out & channel16_Kernel89_Valid_Out & channel17_Kernel89_Valid_Out & channel18_Kernel89_Valid_Out & channel19_Kernel89_Valid_Out & channel20_Kernel89_Valid_Out & channel21_Kernel89_Valid_Out & channel22_Kernel89_Valid_Out & channel23_Kernel89_Valid_Out & channel24_Kernel89_Valid_Out & channel25_Kernel89_Valid_Out & channel26_Kernel89_Valid_Out & channel27_Kernel89_Valid_Out & channel28_Kernel89_Valid_Out & channel29_Kernel89_Valid_Out & channel30_Kernel89_Valid_Out & channel31_Kernel89_Valid_Out & channel32_Kernel89_Valid_Out & channel33_Kernel89_Valid_Out & channel34_Kernel89_Valid_Out & channel35_Kernel89_Valid_Out & channel36_Kernel89_Valid_Out & channel37_Kernel89_Valid_Out & channel38_Kernel89_Valid_Out & channel39_Kernel89_Valid_Out & channel40_Kernel89_Valid_Out & channel41_Kernel89_Valid_Out & channel42_Kernel89_Valid_Out & channel43_Kernel89_Valid_Out & channel44_Kernel89_Valid_Out & channel45_Kernel89_Valid_Out & channel46_Kernel89_Valid_Out & channel47_Kernel89_Valid_Out & channel48_Kernel89_Valid_Out & channel49_Kernel89_Valid_Out & channel50_Kernel89_Valid_Out & channel51_Kernel89_Valid_Out & channel52_Kernel89_Valid_Out & channel53_Kernel89_Valid_Out & channel54_Kernel89_Valid_Out & channel55_Kernel89_Valid_Out & channel56_Kernel89_Valid_Out & channel57_Kernel89_Valid_Out & channel58_Kernel89_Valid_Out & channel59_Kernel89_Valid_Out & channel60_Kernel89_Valid_Out & channel61_Kernel89_Valid_Out & channel62_Kernel89_Valid_Out & channel63_Kernel89_Valid_Out & channel64_Kernel89_Valid_Out;

	wire channel1_Kernel90_Valid_Out, channel2_Kernel90_Valid_Out, channel3_Kernel90_Valid_Out, channel4_Kernel90_Valid_Out, channel5_Kernel90_Valid_Out, channel6_Kernel90_Valid_Out, channel7_Kernel90_Valid_Out, channel8_Kernel90_Valid_Out, channel9_Kernel90_Valid_Out, channel10_Kernel90_Valid_Out, channel11_Kernel90_Valid_Out, channel12_Kernel90_Valid_Out, channel13_Kernel90_Valid_Out, channel14_Kernel90_Valid_Out, channel15_Kernel90_Valid_Out, channel16_Kernel90_Valid_Out, channel17_Kernel90_Valid_Out, channel18_Kernel90_Valid_Out, channel19_Kernel90_Valid_Out, channel20_Kernel90_Valid_Out, channel21_Kernel90_Valid_Out, channel22_Kernel90_Valid_Out, channel23_Kernel90_Valid_Out, channel24_Kernel90_Valid_Out, channel25_Kernel90_Valid_Out, channel26_Kernel90_Valid_Out, channel27_Kernel90_Valid_Out, channel28_Kernel90_Valid_Out, channel29_Kernel90_Valid_Out, channel30_Kernel90_Valid_Out, channel31_Kernel90_Valid_Out, channel32_Kernel90_Valid_Out, channel33_Kernel90_Valid_Out, channel34_Kernel90_Valid_Out, channel35_Kernel90_Valid_Out, channel36_Kernel90_Valid_Out, channel37_Kernel90_Valid_Out, channel38_Kernel90_Valid_Out, channel39_Kernel90_Valid_Out, channel40_Kernel90_Valid_Out, channel41_Kernel90_Valid_Out, channel42_Kernel90_Valid_Out, channel43_Kernel90_Valid_Out, channel44_Kernel90_Valid_Out, channel45_Kernel90_Valid_Out, channel46_Kernel90_Valid_Out, channel47_Kernel90_Valid_Out, channel48_Kernel90_Valid_Out, channel49_Kernel90_Valid_Out, channel50_Kernel90_Valid_Out, channel51_Kernel90_Valid_Out, channel52_Kernel90_Valid_Out, channel53_Kernel90_Valid_Out, channel54_Kernel90_Valid_Out, channel55_Kernel90_Valid_Out, channel56_Kernel90_Valid_Out, channel57_Kernel90_Valid_Out, channel58_Kernel90_Valid_Out, channel59_Kernel90_Valid_Out, channel60_Kernel90_Valid_Out, channel61_Kernel90_Valid_Out, channel62_Kernel90_Valid_Out, channel63_Kernel90_Valid_Out, channel64_Kernel90_Valid_Out;

	assign add_kernel90=channel1_Kernel90_Valid_Out & channel2_Kernel90_Valid_Out & channel3_Kernel90_Valid_Out & channel4_Kernel90_Valid_Out & channel5_Kernel90_Valid_Out & channel6_Kernel90_Valid_Out & channel7_Kernel90_Valid_Out & channel8_Kernel90_Valid_Out & channel9_Kernel90_Valid_Out & channel10_Kernel90_Valid_Out & channel11_Kernel90_Valid_Out & channel12_Kernel90_Valid_Out & channel13_Kernel90_Valid_Out & channel14_Kernel90_Valid_Out & channel15_Kernel90_Valid_Out & channel16_Kernel90_Valid_Out & channel17_Kernel90_Valid_Out & channel18_Kernel90_Valid_Out & channel19_Kernel90_Valid_Out & channel20_Kernel90_Valid_Out & channel21_Kernel90_Valid_Out & channel22_Kernel90_Valid_Out & channel23_Kernel90_Valid_Out & channel24_Kernel90_Valid_Out & channel25_Kernel90_Valid_Out & channel26_Kernel90_Valid_Out & channel27_Kernel90_Valid_Out & channel28_Kernel90_Valid_Out & channel29_Kernel90_Valid_Out & channel30_Kernel90_Valid_Out & channel31_Kernel90_Valid_Out & channel32_Kernel90_Valid_Out & channel33_Kernel90_Valid_Out & channel34_Kernel90_Valid_Out & channel35_Kernel90_Valid_Out & channel36_Kernel90_Valid_Out & channel37_Kernel90_Valid_Out & channel38_Kernel90_Valid_Out & channel39_Kernel90_Valid_Out & channel40_Kernel90_Valid_Out & channel41_Kernel90_Valid_Out & channel42_Kernel90_Valid_Out & channel43_Kernel90_Valid_Out & channel44_Kernel90_Valid_Out & channel45_Kernel90_Valid_Out & channel46_Kernel90_Valid_Out & channel47_Kernel90_Valid_Out & channel48_Kernel90_Valid_Out & channel49_Kernel90_Valid_Out & channel50_Kernel90_Valid_Out & channel51_Kernel90_Valid_Out & channel52_Kernel90_Valid_Out & channel53_Kernel90_Valid_Out & channel54_Kernel90_Valid_Out & channel55_Kernel90_Valid_Out & channel56_Kernel90_Valid_Out & channel57_Kernel90_Valid_Out & channel58_Kernel90_Valid_Out & channel59_Kernel90_Valid_Out & channel60_Kernel90_Valid_Out & channel61_Kernel90_Valid_Out & channel62_Kernel90_Valid_Out & channel63_Kernel90_Valid_Out & channel64_Kernel90_Valid_Out;

	wire channel1_Kernel91_Valid_Out, channel2_Kernel91_Valid_Out, channel3_Kernel91_Valid_Out, channel4_Kernel91_Valid_Out, channel5_Kernel91_Valid_Out, channel6_Kernel91_Valid_Out, channel7_Kernel91_Valid_Out, channel8_Kernel91_Valid_Out, channel9_Kernel91_Valid_Out, channel10_Kernel91_Valid_Out, channel11_Kernel91_Valid_Out, channel12_Kernel91_Valid_Out, channel13_Kernel91_Valid_Out, channel14_Kernel91_Valid_Out, channel15_Kernel91_Valid_Out, channel16_Kernel91_Valid_Out, channel17_Kernel91_Valid_Out, channel18_Kernel91_Valid_Out, channel19_Kernel91_Valid_Out, channel20_Kernel91_Valid_Out, channel21_Kernel91_Valid_Out, channel22_Kernel91_Valid_Out, channel23_Kernel91_Valid_Out, channel24_Kernel91_Valid_Out, channel25_Kernel91_Valid_Out, channel26_Kernel91_Valid_Out, channel27_Kernel91_Valid_Out, channel28_Kernel91_Valid_Out, channel29_Kernel91_Valid_Out, channel30_Kernel91_Valid_Out, channel31_Kernel91_Valid_Out, channel32_Kernel91_Valid_Out, channel33_Kernel91_Valid_Out, channel34_Kernel91_Valid_Out, channel35_Kernel91_Valid_Out, channel36_Kernel91_Valid_Out, channel37_Kernel91_Valid_Out, channel38_Kernel91_Valid_Out, channel39_Kernel91_Valid_Out, channel40_Kernel91_Valid_Out, channel41_Kernel91_Valid_Out, channel42_Kernel91_Valid_Out, channel43_Kernel91_Valid_Out, channel44_Kernel91_Valid_Out, channel45_Kernel91_Valid_Out, channel46_Kernel91_Valid_Out, channel47_Kernel91_Valid_Out, channel48_Kernel91_Valid_Out, channel49_Kernel91_Valid_Out, channel50_Kernel91_Valid_Out, channel51_Kernel91_Valid_Out, channel52_Kernel91_Valid_Out, channel53_Kernel91_Valid_Out, channel54_Kernel91_Valid_Out, channel55_Kernel91_Valid_Out, channel56_Kernel91_Valid_Out, channel57_Kernel91_Valid_Out, channel58_Kernel91_Valid_Out, channel59_Kernel91_Valid_Out, channel60_Kernel91_Valid_Out, channel61_Kernel91_Valid_Out, channel62_Kernel91_Valid_Out, channel63_Kernel91_Valid_Out, channel64_Kernel91_Valid_Out;

	assign add_kernel91=channel1_Kernel91_Valid_Out & channel2_Kernel91_Valid_Out & channel3_Kernel91_Valid_Out & channel4_Kernel91_Valid_Out & channel5_Kernel91_Valid_Out & channel6_Kernel91_Valid_Out & channel7_Kernel91_Valid_Out & channel8_Kernel91_Valid_Out & channel9_Kernel91_Valid_Out & channel10_Kernel91_Valid_Out & channel11_Kernel91_Valid_Out & channel12_Kernel91_Valid_Out & channel13_Kernel91_Valid_Out & channel14_Kernel91_Valid_Out & channel15_Kernel91_Valid_Out & channel16_Kernel91_Valid_Out & channel17_Kernel91_Valid_Out & channel18_Kernel91_Valid_Out & channel19_Kernel91_Valid_Out & channel20_Kernel91_Valid_Out & channel21_Kernel91_Valid_Out & channel22_Kernel91_Valid_Out & channel23_Kernel91_Valid_Out & channel24_Kernel91_Valid_Out & channel25_Kernel91_Valid_Out & channel26_Kernel91_Valid_Out & channel27_Kernel91_Valid_Out & channel28_Kernel91_Valid_Out & channel29_Kernel91_Valid_Out & channel30_Kernel91_Valid_Out & channel31_Kernel91_Valid_Out & channel32_Kernel91_Valid_Out & channel33_Kernel91_Valid_Out & channel34_Kernel91_Valid_Out & channel35_Kernel91_Valid_Out & channel36_Kernel91_Valid_Out & channel37_Kernel91_Valid_Out & channel38_Kernel91_Valid_Out & channel39_Kernel91_Valid_Out & channel40_Kernel91_Valid_Out & channel41_Kernel91_Valid_Out & channel42_Kernel91_Valid_Out & channel43_Kernel91_Valid_Out & channel44_Kernel91_Valid_Out & channel45_Kernel91_Valid_Out & channel46_Kernel91_Valid_Out & channel47_Kernel91_Valid_Out & channel48_Kernel91_Valid_Out & channel49_Kernel91_Valid_Out & channel50_Kernel91_Valid_Out & channel51_Kernel91_Valid_Out & channel52_Kernel91_Valid_Out & channel53_Kernel91_Valid_Out & channel54_Kernel91_Valid_Out & channel55_Kernel91_Valid_Out & channel56_Kernel91_Valid_Out & channel57_Kernel91_Valid_Out & channel58_Kernel91_Valid_Out & channel59_Kernel91_Valid_Out & channel60_Kernel91_Valid_Out & channel61_Kernel91_Valid_Out & channel62_Kernel91_Valid_Out & channel63_Kernel91_Valid_Out & channel64_Kernel91_Valid_Out;

	wire channel1_Kernel92_Valid_Out, channel2_Kernel92_Valid_Out, channel3_Kernel92_Valid_Out, channel4_Kernel92_Valid_Out, channel5_Kernel92_Valid_Out, channel6_Kernel92_Valid_Out, channel7_Kernel92_Valid_Out, channel8_Kernel92_Valid_Out, channel9_Kernel92_Valid_Out, channel10_Kernel92_Valid_Out, channel11_Kernel92_Valid_Out, channel12_Kernel92_Valid_Out, channel13_Kernel92_Valid_Out, channel14_Kernel92_Valid_Out, channel15_Kernel92_Valid_Out, channel16_Kernel92_Valid_Out, channel17_Kernel92_Valid_Out, channel18_Kernel92_Valid_Out, channel19_Kernel92_Valid_Out, channel20_Kernel92_Valid_Out, channel21_Kernel92_Valid_Out, channel22_Kernel92_Valid_Out, channel23_Kernel92_Valid_Out, channel24_Kernel92_Valid_Out, channel25_Kernel92_Valid_Out, channel26_Kernel92_Valid_Out, channel27_Kernel92_Valid_Out, channel28_Kernel92_Valid_Out, channel29_Kernel92_Valid_Out, channel30_Kernel92_Valid_Out, channel31_Kernel92_Valid_Out, channel32_Kernel92_Valid_Out, channel33_Kernel92_Valid_Out, channel34_Kernel92_Valid_Out, channel35_Kernel92_Valid_Out, channel36_Kernel92_Valid_Out, channel37_Kernel92_Valid_Out, channel38_Kernel92_Valid_Out, channel39_Kernel92_Valid_Out, channel40_Kernel92_Valid_Out, channel41_Kernel92_Valid_Out, channel42_Kernel92_Valid_Out, channel43_Kernel92_Valid_Out, channel44_Kernel92_Valid_Out, channel45_Kernel92_Valid_Out, channel46_Kernel92_Valid_Out, channel47_Kernel92_Valid_Out, channel48_Kernel92_Valid_Out, channel49_Kernel92_Valid_Out, channel50_Kernel92_Valid_Out, channel51_Kernel92_Valid_Out, channel52_Kernel92_Valid_Out, channel53_Kernel92_Valid_Out, channel54_Kernel92_Valid_Out, channel55_Kernel92_Valid_Out, channel56_Kernel92_Valid_Out, channel57_Kernel92_Valid_Out, channel58_Kernel92_Valid_Out, channel59_Kernel92_Valid_Out, channel60_Kernel92_Valid_Out, channel61_Kernel92_Valid_Out, channel62_Kernel92_Valid_Out, channel63_Kernel92_Valid_Out, channel64_Kernel92_Valid_Out;

	assign add_kernel92=channel1_Kernel92_Valid_Out & channel2_Kernel92_Valid_Out & channel3_Kernel92_Valid_Out & channel4_Kernel92_Valid_Out & channel5_Kernel92_Valid_Out & channel6_Kernel92_Valid_Out & channel7_Kernel92_Valid_Out & channel8_Kernel92_Valid_Out & channel9_Kernel92_Valid_Out & channel10_Kernel92_Valid_Out & channel11_Kernel92_Valid_Out & channel12_Kernel92_Valid_Out & channel13_Kernel92_Valid_Out & channel14_Kernel92_Valid_Out & channel15_Kernel92_Valid_Out & channel16_Kernel92_Valid_Out & channel17_Kernel92_Valid_Out & channel18_Kernel92_Valid_Out & channel19_Kernel92_Valid_Out & channel20_Kernel92_Valid_Out & channel21_Kernel92_Valid_Out & channel22_Kernel92_Valid_Out & channel23_Kernel92_Valid_Out & channel24_Kernel92_Valid_Out & channel25_Kernel92_Valid_Out & channel26_Kernel92_Valid_Out & channel27_Kernel92_Valid_Out & channel28_Kernel92_Valid_Out & channel29_Kernel92_Valid_Out & channel30_Kernel92_Valid_Out & channel31_Kernel92_Valid_Out & channel32_Kernel92_Valid_Out & channel33_Kernel92_Valid_Out & channel34_Kernel92_Valid_Out & channel35_Kernel92_Valid_Out & channel36_Kernel92_Valid_Out & channel37_Kernel92_Valid_Out & channel38_Kernel92_Valid_Out & channel39_Kernel92_Valid_Out & channel40_Kernel92_Valid_Out & channel41_Kernel92_Valid_Out & channel42_Kernel92_Valid_Out & channel43_Kernel92_Valid_Out & channel44_Kernel92_Valid_Out & channel45_Kernel92_Valid_Out & channel46_Kernel92_Valid_Out & channel47_Kernel92_Valid_Out & channel48_Kernel92_Valid_Out & channel49_Kernel92_Valid_Out & channel50_Kernel92_Valid_Out & channel51_Kernel92_Valid_Out & channel52_Kernel92_Valid_Out & channel53_Kernel92_Valid_Out & channel54_Kernel92_Valid_Out & channel55_Kernel92_Valid_Out & channel56_Kernel92_Valid_Out & channel57_Kernel92_Valid_Out & channel58_Kernel92_Valid_Out & channel59_Kernel92_Valid_Out & channel60_Kernel92_Valid_Out & channel61_Kernel92_Valid_Out & channel62_Kernel92_Valid_Out & channel63_Kernel92_Valid_Out & channel64_Kernel92_Valid_Out;

	wire channel1_Kernel93_Valid_Out, channel2_Kernel93_Valid_Out, channel3_Kernel93_Valid_Out, channel4_Kernel93_Valid_Out, channel5_Kernel93_Valid_Out, channel6_Kernel93_Valid_Out, channel7_Kernel93_Valid_Out, channel8_Kernel93_Valid_Out, channel9_Kernel93_Valid_Out, channel10_Kernel93_Valid_Out, channel11_Kernel93_Valid_Out, channel12_Kernel93_Valid_Out, channel13_Kernel93_Valid_Out, channel14_Kernel93_Valid_Out, channel15_Kernel93_Valid_Out, channel16_Kernel93_Valid_Out, channel17_Kernel93_Valid_Out, channel18_Kernel93_Valid_Out, channel19_Kernel93_Valid_Out, channel20_Kernel93_Valid_Out, channel21_Kernel93_Valid_Out, channel22_Kernel93_Valid_Out, channel23_Kernel93_Valid_Out, channel24_Kernel93_Valid_Out, channel25_Kernel93_Valid_Out, channel26_Kernel93_Valid_Out, channel27_Kernel93_Valid_Out, channel28_Kernel93_Valid_Out, channel29_Kernel93_Valid_Out, channel30_Kernel93_Valid_Out, channel31_Kernel93_Valid_Out, channel32_Kernel93_Valid_Out, channel33_Kernel93_Valid_Out, channel34_Kernel93_Valid_Out, channel35_Kernel93_Valid_Out, channel36_Kernel93_Valid_Out, channel37_Kernel93_Valid_Out, channel38_Kernel93_Valid_Out, channel39_Kernel93_Valid_Out, channel40_Kernel93_Valid_Out, channel41_Kernel93_Valid_Out, channel42_Kernel93_Valid_Out, channel43_Kernel93_Valid_Out, channel44_Kernel93_Valid_Out, channel45_Kernel93_Valid_Out, channel46_Kernel93_Valid_Out, channel47_Kernel93_Valid_Out, channel48_Kernel93_Valid_Out, channel49_Kernel93_Valid_Out, channel50_Kernel93_Valid_Out, channel51_Kernel93_Valid_Out, channel52_Kernel93_Valid_Out, channel53_Kernel93_Valid_Out, channel54_Kernel93_Valid_Out, channel55_Kernel93_Valid_Out, channel56_Kernel93_Valid_Out, channel57_Kernel93_Valid_Out, channel58_Kernel93_Valid_Out, channel59_Kernel93_Valid_Out, channel60_Kernel93_Valid_Out, channel61_Kernel93_Valid_Out, channel62_Kernel93_Valid_Out, channel63_Kernel93_Valid_Out, channel64_Kernel93_Valid_Out;

	assign add_kernel93=channel1_Kernel93_Valid_Out & channel2_Kernel93_Valid_Out & channel3_Kernel93_Valid_Out & channel4_Kernel93_Valid_Out & channel5_Kernel93_Valid_Out & channel6_Kernel93_Valid_Out & channel7_Kernel93_Valid_Out & channel8_Kernel93_Valid_Out & channel9_Kernel93_Valid_Out & channel10_Kernel93_Valid_Out & channel11_Kernel93_Valid_Out & channel12_Kernel93_Valid_Out & channel13_Kernel93_Valid_Out & channel14_Kernel93_Valid_Out & channel15_Kernel93_Valid_Out & channel16_Kernel93_Valid_Out & channel17_Kernel93_Valid_Out & channel18_Kernel93_Valid_Out & channel19_Kernel93_Valid_Out & channel20_Kernel93_Valid_Out & channel21_Kernel93_Valid_Out & channel22_Kernel93_Valid_Out & channel23_Kernel93_Valid_Out & channel24_Kernel93_Valid_Out & channel25_Kernel93_Valid_Out & channel26_Kernel93_Valid_Out & channel27_Kernel93_Valid_Out & channel28_Kernel93_Valid_Out & channel29_Kernel93_Valid_Out & channel30_Kernel93_Valid_Out & channel31_Kernel93_Valid_Out & channel32_Kernel93_Valid_Out & channel33_Kernel93_Valid_Out & channel34_Kernel93_Valid_Out & channel35_Kernel93_Valid_Out & channel36_Kernel93_Valid_Out & channel37_Kernel93_Valid_Out & channel38_Kernel93_Valid_Out & channel39_Kernel93_Valid_Out & channel40_Kernel93_Valid_Out & channel41_Kernel93_Valid_Out & channel42_Kernel93_Valid_Out & channel43_Kernel93_Valid_Out & channel44_Kernel93_Valid_Out & channel45_Kernel93_Valid_Out & channel46_Kernel93_Valid_Out & channel47_Kernel93_Valid_Out & channel48_Kernel93_Valid_Out & channel49_Kernel93_Valid_Out & channel50_Kernel93_Valid_Out & channel51_Kernel93_Valid_Out & channel52_Kernel93_Valid_Out & channel53_Kernel93_Valid_Out & channel54_Kernel93_Valid_Out & channel55_Kernel93_Valid_Out & channel56_Kernel93_Valid_Out & channel57_Kernel93_Valid_Out & channel58_Kernel93_Valid_Out & channel59_Kernel93_Valid_Out & channel60_Kernel93_Valid_Out & channel61_Kernel93_Valid_Out & channel62_Kernel93_Valid_Out & channel63_Kernel93_Valid_Out & channel64_Kernel93_Valid_Out;

	wire channel1_Kernel94_Valid_Out, channel2_Kernel94_Valid_Out, channel3_Kernel94_Valid_Out, channel4_Kernel94_Valid_Out, channel5_Kernel94_Valid_Out, channel6_Kernel94_Valid_Out, channel7_Kernel94_Valid_Out, channel8_Kernel94_Valid_Out, channel9_Kernel94_Valid_Out, channel10_Kernel94_Valid_Out, channel11_Kernel94_Valid_Out, channel12_Kernel94_Valid_Out, channel13_Kernel94_Valid_Out, channel14_Kernel94_Valid_Out, channel15_Kernel94_Valid_Out, channel16_Kernel94_Valid_Out, channel17_Kernel94_Valid_Out, channel18_Kernel94_Valid_Out, channel19_Kernel94_Valid_Out, channel20_Kernel94_Valid_Out, channel21_Kernel94_Valid_Out, channel22_Kernel94_Valid_Out, channel23_Kernel94_Valid_Out, channel24_Kernel94_Valid_Out, channel25_Kernel94_Valid_Out, channel26_Kernel94_Valid_Out, channel27_Kernel94_Valid_Out, channel28_Kernel94_Valid_Out, channel29_Kernel94_Valid_Out, channel30_Kernel94_Valid_Out, channel31_Kernel94_Valid_Out, channel32_Kernel94_Valid_Out, channel33_Kernel94_Valid_Out, channel34_Kernel94_Valid_Out, channel35_Kernel94_Valid_Out, channel36_Kernel94_Valid_Out, channel37_Kernel94_Valid_Out, channel38_Kernel94_Valid_Out, channel39_Kernel94_Valid_Out, channel40_Kernel94_Valid_Out, channel41_Kernel94_Valid_Out, channel42_Kernel94_Valid_Out, channel43_Kernel94_Valid_Out, channel44_Kernel94_Valid_Out, channel45_Kernel94_Valid_Out, channel46_Kernel94_Valid_Out, channel47_Kernel94_Valid_Out, channel48_Kernel94_Valid_Out, channel49_Kernel94_Valid_Out, channel50_Kernel94_Valid_Out, channel51_Kernel94_Valid_Out, channel52_Kernel94_Valid_Out, channel53_Kernel94_Valid_Out, channel54_Kernel94_Valid_Out, channel55_Kernel94_Valid_Out, channel56_Kernel94_Valid_Out, channel57_Kernel94_Valid_Out, channel58_Kernel94_Valid_Out, channel59_Kernel94_Valid_Out, channel60_Kernel94_Valid_Out, channel61_Kernel94_Valid_Out, channel62_Kernel94_Valid_Out, channel63_Kernel94_Valid_Out, channel64_Kernel94_Valid_Out;

	assign add_kernel94=channel1_Kernel94_Valid_Out & channel2_Kernel94_Valid_Out & channel3_Kernel94_Valid_Out & channel4_Kernel94_Valid_Out & channel5_Kernel94_Valid_Out & channel6_Kernel94_Valid_Out & channel7_Kernel94_Valid_Out & channel8_Kernel94_Valid_Out & channel9_Kernel94_Valid_Out & channel10_Kernel94_Valid_Out & channel11_Kernel94_Valid_Out & channel12_Kernel94_Valid_Out & channel13_Kernel94_Valid_Out & channel14_Kernel94_Valid_Out & channel15_Kernel94_Valid_Out & channel16_Kernel94_Valid_Out & channel17_Kernel94_Valid_Out & channel18_Kernel94_Valid_Out & channel19_Kernel94_Valid_Out & channel20_Kernel94_Valid_Out & channel21_Kernel94_Valid_Out & channel22_Kernel94_Valid_Out & channel23_Kernel94_Valid_Out & channel24_Kernel94_Valid_Out & channel25_Kernel94_Valid_Out & channel26_Kernel94_Valid_Out & channel27_Kernel94_Valid_Out & channel28_Kernel94_Valid_Out & channel29_Kernel94_Valid_Out & channel30_Kernel94_Valid_Out & channel31_Kernel94_Valid_Out & channel32_Kernel94_Valid_Out & channel33_Kernel94_Valid_Out & channel34_Kernel94_Valid_Out & channel35_Kernel94_Valid_Out & channel36_Kernel94_Valid_Out & channel37_Kernel94_Valid_Out & channel38_Kernel94_Valid_Out & channel39_Kernel94_Valid_Out & channel40_Kernel94_Valid_Out & channel41_Kernel94_Valid_Out & channel42_Kernel94_Valid_Out & channel43_Kernel94_Valid_Out & channel44_Kernel94_Valid_Out & channel45_Kernel94_Valid_Out & channel46_Kernel94_Valid_Out & channel47_Kernel94_Valid_Out & channel48_Kernel94_Valid_Out & channel49_Kernel94_Valid_Out & channel50_Kernel94_Valid_Out & channel51_Kernel94_Valid_Out & channel52_Kernel94_Valid_Out & channel53_Kernel94_Valid_Out & channel54_Kernel94_Valid_Out & channel55_Kernel94_Valid_Out & channel56_Kernel94_Valid_Out & channel57_Kernel94_Valid_Out & channel58_Kernel94_Valid_Out & channel59_Kernel94_Valid_Out & channel60_Kernel94_Valid_Out & channel61_Kernel94_Valid_Out & channel62_Kernel94_Valid_Out & channel63_Kernel94_Valid_Out & channel64_Kernel94_Valid_Out;

	wire channel1_Kernel95_Valid_Out, channel2_Kernel95_Valid_Out, channel3_Kernel95_Valid_Out, channel4_Kernel95_Valid_Out, channel5_Kernel95_Valid_Out, channel6_Kernel95_Valid_Out, channel7_Kernel95_Valid_Out, channel8_Kernel95_Valid_Out, channel9_Kernel95_Valid_Out, channel10_Kernel95_Valid_Out, channel11_Kernel95_Valid_Out, channel12_Kernel95_Valid_Out, channel13_Kernel95_Valid_Out, channel14_Kernel95_Valid_Out, channel15_Kernel95_Valid_Out, channel16_Kernel95_Valid_Out, channel17_Kernel95_Valid_Out, channel18_Kernel95_Valid_Out, channel19_Kernel95_Valid_Out, channel20_Kernel95_Valid_Out, channel21_Kernel95_Valid_Out, channel22_Kernel95_Valid_Out, channel23_Kernel95_Valid_Out, channel24_Kernel95_Valid_Out, channel25_Kernel95_Valid_Out, channel26_Kernel95_Valid_Out, channel27_Kernel95_Valid_Out, channel28_Kernel95_Valid_Out, channel29_Kernel95_Valid_Out, channel30_Kernel95_Valid_Out, channel31_Kernel95_Valid_Out, channel32_Kernel95_Valid_Out, channel33_Kernel95_Valid_Out, channel34_Kernel95_Valid_Out, channel35_Kernel95_Valid_Out, channel36_Kernel95_Valid_Out, channel37_Kernel95_Valid_Out, channel38_Kernel95_Valid_Out, channel39_Kernel95_Valid_Out, channel40_Kernel95_Valid_Out, channel41_Kernel95_Valid_Out, channel42_Kernel95_Valid_Out, channel43_Kernel95_Valid_Out, channel44_Kernel95_Valid_Out, channel45_Kernel95_Valid_Out, channel46_Kernel95_Valid_Out, channel47_Kernel95_Valid_Out, channel48_Kernel95_Valid_Out, channel49_Kernel95_Valid_Out, channel50_Kernel95_Valid_Out, channel51_Kernel95_Valid_Out, channel52_Kernel95_Valid_Out, channel53_Kernel95_Valid_Out, channel54_Kernel95_Valid_Out, channel55_Kernel95_Valid_Out, channel56_Kernel95_Valid_Out, channel57_Kernel95_Valid_Out, channel58_Kernel95_Valid_Out, channel59_Kernel95_Valid_Out, channel60_Kernel95_Valid_Out, channel61_Kernel95_Valid_Out, channel62_Kernel95_Valid_Out, channel63_Kernel95_Valid_Out, channel64_Kernel95_Valid_Out;

	assign add_kernel95=channel1_Kernel95_Valid_Out & channel2_Kernel95_Valid_Out & channel3_Kernel95_Valid_Out & channel4_Kernel95_Valid_Out & channel5_Kernel95_Valid_Out & channel6_Kernel95_Valid_Out & channel7_Kernel95_Valid_Out & channel8_Kernel95_Valid_Out & channel9_Kernel95_Valid_Out & channel10_Kernel95_Valid_Out & channel11_Kernel95_Valid_Out & channel12_Kernel95_Valid_Out & channel13_Kernel95_Valid_Out & channel14_Kernel95_Valid_Out & channel15_Kernel95_Valid_Out & channel16_Kernel95_Valid_Out & channel17_Kernel95_Valid_Out & channel18_Kernel95_Valid_Out & channel19_Kernel95_Valid_Out & channel20_Kernel95_Valid_Out & channel21_Kernel95_Valid_Out & channel22_Kernel95_Valid_Out & channel23_Kernel95_Valid_Out & channel24_Kernel95_Valid_Out & channel25_Kernel95_Valid_Out & channel26_Kernel95_Valid_Out & channel27_Kernel95_Valid_Out & channel28_Kernel95_Valid_Out & channel29_Kernel95_Valid_Out & channel30_Kernel95_Valid_Out & channel31_Kernel95_Valid_Out & channel32_Kernel95_Valid_Out & channel33_Kernel95_Valid_Out & channel34_Kernel95_Valid_Out & channel35_Kernel95_Valid_Out & channel36_Kernel95_Valid_Out & channel37_Kernel95_Valid_Out & channel38_Kernel95_Valid_Out & channel39_Kernel95_Valid_Out & channel40_Kernel95_Valid_Out & channel41_Kernel95_Valid_Out & channel42_Kernel95_Valid_Out & channel43_Kernel95_Valid_Out & channel44_Kernel95_Valid_Out & channel45_Kernel95_Valid_Out & channel46_Kernel95_Valid_Out & channel47_Kernel95_Valid_Out & channel48_Kernel95_Valid_Out & channel49_Kernel95_Valid_Out & channel50_Kernel95_Valid_Out & channel51_Kernel95_Valid_Out & channel52_Kernel95_Valid_Out & channel53_Kernel95_Valid_Out & channel54_Kernel95_Valid_Out & channel55_Kernel95_Valid_Out & channel56_Kernel95_Valid_Out & channel57_Kernel95_Valid_Out & channel58_Kernel95_Valid_Out & channel59_Kernel95_Valid_Out & channel60_Kernel95_Valid_Out & channel61_Kernel95_Valid_Out & channel62_Kernel95_Valid_Out & channel63_Kernel95_Valid_Out & channel64_Kernel95_Valid_Out;

	wire channel1_Kernel96_Valid_Out, channel2_Kernel96_Valid_Out, channel3_Kernel96_Valid_Out, channel4_Kernel96_Valid_Out, channel5_Kernel96_Valid_Out, channel6_Kernel96_Valid_Out, channel7_Kernel96_Valid_Out, channel8_Kernel96_Valid_Out, channel9_Kernel96_Valid_Out, channel10_Kernel96_Valid_Out, channel11_Kernel96_Valid_Out, channel12_Kernel96_Valid_Out, channel13_Kernel96_Valid_Out, channel14_Kernel96_Valid_Out, channel15_Kernel96_Valid_Out, channel16_Kernel96_Valid_Out, channel17_Kernel96_Valid_Out, channel18_Kernel96_Valid_Out, channel19_Kernel96_Valid_Out, channel20_Kernel96_Valid_Out, channel21_Kernel96_Valid_Out, channel22_Kernel96_Valid_Out, channel23_Kernel96_Valid_Out, channel24_Kernel96_Valid_Out, channel25_Kernel96_Valid_Out, channel26_Kernel96_Valid_Out, channel27_Kernel96_Valid_Out, channel28_Kernel96_Valid_Out, channel29_Kernel96_Valid_Out, channel30_Kernel96_Valid_Out, channel31_Kernel96_Valid_Out, channel32_Kernel96_Valid_Out, channel33_Kernel96_Valid_Out, channel34_Kernel96_Valid_Out, channel35_Kernel96_Valid_Out, channel36_Kernel96_Valid_Out, channel37_Kernel96_Valid_Out, channel38_Kernel96_Valid_Out, channel39_Kernel96_Valid_Out, channel40_Kernel96_Valid_Out, channel41_Kernel96_Valid_Out, channel42_Kernel96_Valid_Out, channel43_Kernel96_Valid_Out, channel44_Kernel96_Valid_Out, channel45_Kernel96_Valid_Out, channel46_Kernel96_Valid_Out, channel47_Kernel96_Valid_Out, channel48_Kernel96_Valid_Out, channel49_Kernel96_Valid_Out, channel50_Kernel96_Valid_Out, channel51_Kernel96_Valid_Out, channel52_Kernel96_Valid_Out, channel53_Kernel96_Valid_Out, channel54_Kernel96_Valid_Out, channel55_Kernel96_Valid_Out, channel56_Kernel96_Valid_Out, channel57_Kernel96_Valid_Out, channel58_Kernel96_Valid_Out, channel59_Kernel96_Valid_Out, channel60_Kernel96_Valid_Out, channel61_Kernel96_Valid_Out, channel62_Kernel96_Valid_Out, channel63_Kernel96_Valid_Out, channel64_Kernel96_Valid_Out;

	assign add_kernel96=channel1_Kernel96_Valid_Out & channel2_Kernel96_Valid_Out & channel3_Kernel96_Valid_Out & channel4_Kernel96_Valid_Out & channel5_Kernel96_Valid_Out & channel6_Kernel96_Valid_Out & channel7_Kernel96_Valid_Out & channel8_Kernel96_Valid_Out & channel9_Kernel96_Valid_Out & channel10_Kernel96_Valid_Out & channel11_Kernel96_Valid_Out & channel12_Kernel96_Valid_Out & channel13_Kernel96_Valid_Out & channel14_Kernel96_Valid_Out & channel15_Kernel96_Valid_Out & channel16_Kernel96_Valid_Out & channel17_Kernel96_Valid_Out & channel18_Kernel96_Valid_Out & channel19_Kernel96_Valid_Out & channel20_Kernel96_Valid_Out & channel21_Kernel96_Valid_Out & channel22_Kernel96_Valid_Out & channel23_Kernel96_Valid_Out & channel24_Kernel96_Valid_Out & channel25_Kernel96_Valid_Out & channel26_Kernel96_Valid_Out & channel27_Kernel96_Valid_Out & channel28_Kernel96_Valid_Out & channel29_Kernel96_Valid_Out & channel30_Kernel96_Valid_Out & channel31_Kernel96_Valid_Out & channel32_Kernel96_Valid_Out & channel33_Kernel96_Valid_Out & channel34_Kernel96_Valid_Out & channel35_Kernel96_Valid_Out & channel36_Kernel96_Valid_Out & channel37_Kernel96_Valid_Out & channel38_Kernel96_Valid_Out & channel39_Kernel96_Valid_Out & channel40_Kernel96_Valid_Out & channel41_Kernel96_Valid_Out & channel42_Kernel96_Valid_Out & channel43_Kernel96_Valid_Out & channel44_Kernel96_Valid_Out & channel45_Kernel96_Valid_Out & channel46_Kernel96_Valid_Out & channel47_Kernel96_Valid_Out & channel48_Kernel96_Valid_Out & channel49_Kernel96_Valid_Out & channel50_Kernel96_Valid_Out & channel51_Kernel96_Valid_Out & channel52_Kernel96_Valid_Out & channel53_Kernel96_Valid_Out & channel54_Kernel96_Valid_Out & channel55_Kernel96_Valid_Out & channel56_Kernel96_Valid_Out & channel57_Kernel96_Valid_Out & channel58_Kernel96_Valid_Out & channel59_Kernel96_Valid_Out & channel60_Kernel96_Valid_Out & channel61_Kernel96_Valid_Out & channel62_Kernel96_Valid_Out & channel63_Kernel96_Valid_Out & channel64_Kernel96_Valid_Out;

	wire channel1_Kernel97_Valid_Out, channel2_Kernel97_Valid_Out, channel3_Kernel97_Valid_Out, channel4_Kernel97_Valid_Out, channel5_Kernel97_Valid_Out, channel6_Kernel97_Valid_Out, channel7_Kernel97_Valid_Out, channel8_Kernel97_Valid_Out, channel9_Kernel97_Valid_Out, channel10_Kernel97_Valid_Out, channel11_Kernel97_Valid_Out, channel12_Kernel97_Valid_Out, channel13_Kernel97_Valid_Out, channel14_Kernel97_Valid_Out, channel15_Kernel97_Valid_Out, channel16_Kernel97_Valid_Out, channel17_Kernel97_Valid_Out, channel18_Kernel97_Valid_Out, channel19_Kernel97_Valid_Out, channel20_Kernel97_Valid_Out, channel21_Kernel97_Valid_Out, channel22_Kernel97_Valid_Out, channel23_Kernel97_Valid_Out, channel24_Kernel97_Valid_Out, channel25_Kernel97_Valid_Out, channel26_Kernel97_Valid_Out, channel27_Kernel97_Valid_Out, channel28_Kernel97_Valid_Out, channel29_Kernel97_Valid_Out, channel30_Kernel97_Valid_Out, channel31_Kernel97_Valid_Out, channel32_Kernel97_Valid_Out, channel33_Kernel97_Valid_Out, channel34_Kernel97_Valid_Out, channel35_Kernel97_Valid_Out, channel36_Kernel97_Valid_Out, channel37_Kernel97_Valid_Out, channel38_Kernel97_Valid_Out, channel39_Kernel97_Valid_Out, channel40_Kernel97_Valid_Out, channel41_Kernel97_Valid_Out, channel42_Kernel97_Valid_Out, channel43_Kernel97_Valid_Out, channel44_Kernel97_Valid_Out, channel45_Kernel97_Valid_Out, channel46_Kernel97_Valid_Out, channel47_Kernel97_Valid_Out, channel48_Kernel97_Valid_Out, channel49_Kernel97_Valid_Out, channel50_Kernel97_Valid_Out, channel51_Kernel97_Valid_Out, channel52_Kernel97_Valid_Out, channel53_Kernel97_Valid_Out, channel54_Kernel97_Valid_Out, channel55_Kernel97_Valid_Out, channel56_Kernel97_Valid_Out, channel57_Kernel97_Valid_Out, channel58_Kernel97_Valid_Out, channel59_Kernel97_Valid_Out, channel60_Kernel97_Valid_Out, channel61_Kernel97_Valid_Out, channel62_Kernel97_Valid_Out, channel63_Kernel97_Valid_Out, channel64_Kernel97_Valid_Out;

	assign add_kernel97=channel1_Kernel97_Valid_Out & channel2_Kernel97_Valid_Out & channel3_Kernel97_Valid_Out & channel4_Kernel97_Valid_Out & channel5_Kernel97_Valid_Out & channel6_Kernel97_Valid_Out & channel7_Kernel97_Valid_Out & channel8_Kernel97_Valid_Out & channel9_Kernel97_Valid_Out & channel10_Kernel97_Valid_Out & channel11_Kernel97_Valid_Out & channel12_Kernel97_Valid_Out & channel13_Kernel97_Valid_Out & channel14_Kernel97_Valid_Out & channel15_Kernel97_Valid_Out & channel16_Kernel97_Valid_Out & channel17_Kernel97_Valid_Out & channel18_Kernel97_Valid_Out & channel19_Kernel97_Valid_Out & channel20_Kernel97_Valid_Out & channel21_Kernel97_Valid_Out & channel22_Kernel97_Valid_Out & channel23_Kernel97_Valid_Out & channel24_Kernel97_Valid_Out & channel25_Kernel97_Valid_Out & channel26_Kernel97_Valid_Out & channel27_Kernel97_Valid_Out & channel28_Kernel97_Valid_Out & channel29_Kernel97_Valid_Out & channel30_Kernel97_Valid_Out & channel31_Kernel97_Valid_Out & channel32_Kernel97_Valid_Out & channel33_Kernel97_Valid_Out & channel34_Kernel97_Valid_Out & channel35_Kernel97_Valid_Out & channel36_Kernel97_Valid_Out & channel37_Kernel97_Valid_Out & channel38_Kernel97_Valid_Out & channel39_Kernel97_Valid_Out & channel40_Kernel97_Valid_Out & channel41_Kernel97_Valid_Out & channel42_Kernel97_Valid_Out & channel43_Kernel97_Valid_Out & channel44_Kernel97_Valid_Out & channel45_Kernel97_Valid_Out & channel46_Kernel97_Valid_Out & channel47_Kernel97_Valid_Out & channel48_Kernel97_Valid_Out & channel49_Kernel97_Valid_Out & channel50_Kernel97_Valid_Out & channel51_Kernel97_Valid_Out & channel52_Kernel97_Valid_Out & channel53_Kernel97_Valid_Out & channel54_Kernel97_Valid_Out & channel55_Kernel97_Valid_Out & channel56_Kernel97_Valid_Out & channel57_Kernel97_Valid_Out & channel58_Kernel97_Valid_Out & channel59_Kernel97_Valid_Out & channel60_Kernel97_Valid_Out & channel61_Kernel97_Valid_Out & channel62_Kernel97_Valid_Out & channel63_Kernel97_Valid_Out & channel64_Kernel97_Valid_Out;

	wire channel1_Kernel98_Valid_Out, channel2_Kernel98_Valid_Out, channel3_Kernel98_Valid_Out, channel4_Kernel98_Valid_Out, channel5_Kernel98_Valid_Out, channel6_Kernel98_Valid_Out, channel7_Kernel98_Valid_Out, channel8_Kernel98_Valid_Out, channel9_Kernel98_Valid_Out, channel10_Kernel98_Valid_Out, channel11_Kernel98_Valid_Out, channel12_Kernel98_Valid_Out, channel13_Kernel98_Valid_Out, channel14_Kernel98_Valid_Out, channel15_Kernel98_Valid_Out, channel16_Kernel98_Valid_Out, channel17_Kernel98_Valid_Out, channel18_Kernel98_Valid_Out, channel19_Kernel98_Valid_Out, channel20_Kernel98_Valid_Out, channel21_Kernel98_Valid_Out, channel22_Kernel98_Valid_Out, channel23_Kernel98_Valid_Out, channel24_Kernel98_Valid_Out, channel25_Kernel98_Valid_Out, channel26_Kernel98_Valid_Out, channel27_Kernel98_Valid_Out, channel28_Kernel98_Valid_Out, channel29_Kernel98_Valid_Out, channel30_Kernel98_Valid_Out, channel31_Kernel98_Valid_Out, channel32_Kernel98_Valid_Out, channel33_Kernel98_Valid_Out, channel34_Kernel98_Valid_Out, channel35_Kernel98_Valid_Out, channel36_Kernel98_Valid_Out, channel37_Kernel98_Valid_Out, channel38_Kernel98_Valid_Out, channel39_Kernel98_Valid_Out, channel40_Kernel98_Valid_Out, channel41_Kernel98_Valid_Out, channel42_Kernel98_Valid_Out, channel43_Kernel98_Valid_Out, channel44_Kernel98_Valid_Out, channel45_Kernel98_Valid_Out, channel46_Kernel98_Valid_Out, channel47_Kernel98_Valid_Out, channel48_Kernel98_Valid_Out, channel49_Kernel98_Valid_Out, channel50_Kernel98_Valid_Out, channel51_Kernel98_Valid_Out, channel52_Kernel98_Valid_Out, channel53_Kernel98_Valid_Out, channel54_Kernel98_Valid_Out, channel55_Kernel98_Valid_Out, channel56_Kernel98_Valid_Out, channel57_Kernel98_Valid_Out, channel58_Kernel98_Valid_Out, channel59_Kernel98_Valid_Out, channel60_Kernel98_Valid_Out, channel61_Kernel98_Valid_Out, channel62_Kernel98_Valid_Out, channel63_Kernel98_Valid_Out, channel64_Kernel98_Valid_Out;

	assign add_kernel98=channel1_Kernel98_Valid_Out & channel2_Kernel98_Valid_Out & channel3_Kernel98_Valid_Out & channel4_Kernel98_Valid_Out & channel5_Kernel98_Valid_Out & channel6_Kernel98_Valid_Out & channel7_Kernel98_Valid_Out & channel8_Kernel98_Valid_Out & channel9_Kernel98_Valid_Out & channel10_Kernel98_Valid_Out & channel11_Kernel98_Valid_Out & channel12_Kernel98_Valid_Out & channel13_Kernel98_Valid_Out & channel14_Kernel98_Valid_Out & channel15_Kernel98_Valid_Out & channel16_Kernel98_Valid_Out & channel17_Kernel98_Valid_Out & channel18_Kernel98_Valid_Out & channel19_Kernel98_Valid_Out & channel20_Kernel98_Valid_Out & channel21_Kernel98_Valid_Out & channel22_Kernel98_Valid_Out & channel23_Kernel98_Valid_Out & channel24_Kernel98_Valid_Out & channel25_Kernel98_Valid_Out & channel26_Kernel98_Valid_Out & channel27_Kernel98_Valid_Out & channel28_Kernel98_Valid_Out & channel29_Kernel98_Valid_Out & channel30_Kernel98_Valid_Out & channel31_Kernel98_Valid_Out & channel32_Kernel98_Valid_Out & channel33_Kernel98_Valid_Out & channel34_Kernel98_Valid_Out & channel35_Kernel98_Valid_Out & channel36_Kernel98_Valid_Out & channel37_Kernel98_Valid_Out & channel38_Kernel98_Valid_Out & channel39_Kernel98_Valid_Out & channel40_Kernel98_Valid_Out & channel41_Kernel98_Valid_Out & channel42_Kernel98_Valid_Out & channel43_Kernel98_Valid_Out & channel44_Kernel98_Valid_Out & channel45_Kernel98_Valid_Out & channel46_Kernel98_Valid_Out & channel47_Kernel98_Valid_Out & channel48_Kernel98_Valid_Out & channel49_Kernel98_Valid_Out & channel50_Kernel98_Valid_Out & channel51_Kernel98_Valid_Out & channel52_Kernel98_Valid_Out & channel53_Kernel98_Valid_Out & channel54_Kernel98_Valid_Out & channel55_Kernel98_Valid_Out & channel56_Kernel98_Valid_Out & channel57_Kernel98_Valid_Out & channel58_Kernel98_Valid_Out & channel59_Kernel98_Valid_Out & channel60_Kernel98_Valid_Out & channel61_Kernel98_Valid_Out & channel62_Kernel98_Valid_Out & channel63_Kernel98_Valid_Out & channel64_Kernel98_Valid_Out;

	wire channel1_Kernel99_Valid_Out, channel2_Kernel99_Valid_Out, channel3_Kernel99_Valid_Out, channel4_Kernel99_Valid_Out, channel5_Kernel99_Valid_Out, channel6_Kernel99_Valid_Out, channel7_Kernel99_Valid_Out, channel8_Kernel99_Valid_Out, channel9_Kernel99_Valid_Out, channel10_Kernel99_Valid_Out, channel11_Kernel99_Valid_Out, channel12_Kernel99_Valid_Out, channel13_Kernel99_Valid_Out, channel14_Kernel99_Valid_Out, channel15_Kernel99_Valid_Out, channel16_Kernel99_Valid_Out, channel17_Kernel99_Valid_Out, channel18_Kernel99_Valid_Out, channel19_Kernel99_Valid_Out, channel20_Kernel99_Valid_Out, channel21_Kernel99_Valid_Out, channel22_Kernel99_Valid_Out, channel23_Kernel99_Valid_Out, channel24_Kernel99_Valid_Out, channel25_Kernel99_Valid_Out, channel26_Kernel99_Valid_Out, channel27_Kernel99_Valid_Out, channel28_Kernel99_Valid_Out, channel29_Kernel99_Valid_Out, channel30_Kernel99_Valid_Out, channel31_Kernel99_Valid_Out, channel32_Kernel99_Valid_Out, channel33_Kernel99_Valid_Out, channel34_Kernel99_Valid_Out, channel35_Kernel99_Valid_Out, channel36_Kernel99_Valid_Out, channel37_Kernel99_Valid_Out, channel38_Kernel99_Valid_Out, channel39_Kernel99_Valid_Out, channel40_Kernel99_Valid_Out, channel41_Kernel99_Valid_Out, channel42_Kernel99_Valid_Out, channel43_Kernel99_Valid_Out, channel44_Kernel99_Valid_Out, channel45_Kernel99_Valid_Out, channel46_Kernel99_Valid_Out, channel47_Kernel99_Valid_Out, channel48_Kernel99_Valid_Out, channel49_Kernel99_Valid_Out, channel50_Kernel99_Valid_Out, channel51_Kernel99_Valid_Out, channel52_Kernel99_Valid_Out, channel53_Kernel99_Valid_Out, channel54_Kernel99_Valid_Out, channel55_Kernel99_Valid_Out, channel56_Kernel99_Valid_Out, channel57_Kernel99_Valid_Out, channel58_Kernel99_Valid_Out, channel59_Kernel99_Valid_Out, channel60_Kernel99_Valid_Out, channel61_Kernel99_Valid_Out, channel62_Kernel99_Valid_Out, channel63_Kernel99_Valid_Out, channel64_Kernel99_Valid_Out;

	assign add_kernel99=channel1_Kernel99_Valid_Out & channel2_Kernel99_Valid_Out & channel3_Kernel99_Valid_Out & channel4_Kernel99_Valid_Out & channel5_Kernel99_Valid_Out & channel6_Kernel99_Valid_Out & channel7_Kernel99_Valid_Out & channel8_Kernel99_Valid_Out & channel9_Kernel99_Valid_Out & channel10_Kernel99_Valid_Out & channel11_Kernel99_Valid_Out & channel12_Kernel99_Valid_Out & channel13_Kernel99_Valid_Out & channel14_Kernel99_Valid_Out & channel15_Kernel99_Valid_Out & channel16_Kernel99_Valid_Out & channel17_Kernel99_Valid_Out & channel18_Kernel99_Valid_Out & channel19_Kernel99_Valid_Out & channel20_Kernel99_Valid_Out & channel21_Kernel99_Valid_Out & channel22_Kernel99_Valid_Out & channel23_Kernel99_Valid_Out & channel24_Kernel99_Valid_Out & channel25_Kernel99_Valid_Out & channel26_Kernel99_Valid_Out & channel27_Kernel99_Valid_Out & channel28_Kernel99_Valid_Out & channel29_Kernel99_Valid_Out & channel30_Kernel99_Valid_Out & channel31_Kernel99_Valid_Out & channel32_Kernel99_Valid_Out & channel33_Kernel99_Valid_Out & channel34_Kernel99_Valid_Out & channel35_Kernel99_Valid_Out & channel36_Kernel99_Valid_Out & channel37_Kernel99_Valid_Out & channel38_Kernel99_Valid_Out & channel39_Kernel99_Valid_Out & channel40_Kernel99_Valid_Out & channel41_Kernel99_Valid_Out & channel42_Kernel99_Valid_Out & channel43_Kernel99_Valid_Out & channel44_Kernel99_Valid_Out & channel45_Kernel99_Valid_Out & channel46_Kernel99_Valid_Out & channel47_Kernel99_Valid_Out & channel48_Kernel99_Valid_Out & channel49_Kernel99_Valid_Out & channel50_Kernel99_Valid_Out & channel51_Kernel99_Valid_Out & channel52_Kernel99_Valid_Out & channel53_Kernel99_Valid_Out & channel54_Kernel99_Valid_Out & channel55_Kernel99_Valid_Out & channel56_Kernel99_Valid_Out & channel57_Kernel99_Valid_Out & channel58_Kernel99_Valid_Out & channel59_Kernel99_Valid_Out & channel60_Kernel99_Valid_Out & channel61_Kernel99_Valid_Out & channel62_Kernel99_Valid_Out & channel63_Kernel99_Valid_Out & channel64_Kernel99_Valid_Out;

	wire channel1_Kernel100_Valid_Out, channel2_Kernel100_Valid_Out, channel3_Kernel100_Valid_Out, channel4_Kernel100_Valid_Out, channel5_Kernel100_Valid_Out, channel6_Kernel100_Valid_Out, channel7_Kernel100_Valid_Out, channel8_Kernel100_Valid_Out, channel9_Kernel100_Valid_Out, channel10_Kernel100_Valid_Out, channel11_Kernel100_Valid_Out, channel12_Kernel100_Valid_Out, channel13_Kernel100_Valid_Out, channel14_Kernel100_Valid_Out, channel15_Kernel100_Valid_Out, channel16_Kernel100_Valid_Out, channel17_Kernel100_Valid_Out, channel18_Kernel100_Valid_Out, channel19_Kernel100_Valid_Out, channel20_Kernel100_Valid_Out, channel21_Kernel100_Valid_Out, channel22_Kernel100_Valid_Out, channel23_Kernel100_Valid_Out, channel24_Kernel100_Valid_Out, channel25_Kernel100_Valid_Out, channel26_Kernel100_Valid_Out, channel27_Kernel100_Valid_Out, channel28_Kernel100_Valid_Out, channel29_Kernel100_Valid_Out, channel30_Kernel100_Valid_Out, channel31_Kernel100_Valid_Out, channel32_Kernel100_Valid_Out, channel33_Kernel100_Valid_Out, channel34_Kernel100_Valid_Out, channel35_Kernel100_Valid_Out, channel36_Kernel100_Valid_Out, channel37_Kernel100_Valid_Out, channel38_Kernel100_Valid_Out, channel39_Kernel100_Valid_Out, channel40_Kernel100_Valid_Out, channel41_Kernel100_Valid_Out, channel42_Kernel100_Valid_Out, channel43_Kernel100_Valid_Out, channel44_Kernel100_Valid_Out, channel45_Kernel100_Valid_Out, channel46_Kernel100_Valid_Out, channel47_Kernel100_Valid_Out, channel48_Kernel100_Valid_Out, channel49_Kernel100_Valid_Out, channel50_Kernel100_Valid_Out, channel51_Kernel100_Valid_Out, channel52_Kernel100_Valid_Out, channel53_Kernel100_Valid_Out, channel54_Kernel100_Valid_Out, channel55_Kernel100_Valid_Out, channel56_Kernel100_Valid_Out, channel57_Kernel100_Valid_Out, channel58_Kernel100_Valid_Out, channel59_Kernel100_Valid_Out, channel60_Kernel100_Valid_Out, channel61_Kernel100_Valid_Out, channel62_Kernel100_Valid_Out, channel63_Kernel100_Valid_Out, channel64_Kernel100_Valid_Out;

	assign add_kernel100=channel1_Kernel100_Valid_Out & channel2_Kernel100_Valid_Out & channel3_Kernel100_Valid_Out & channel4_Kernel100_Valid_Out & channel5_Kernel100_Valid_Out & channel6_Kernel100_Valid_Out & channel7_Kernel100_Valid_Out & channel8_Kernel100_Valid_Out & channel9_Kernel100_Valid_Out & channel10_Kernel100_Valid_Out & channel11_Kernel100_Valid_Out & channel12_Kernel100_Valid_Out & channel13_Kernel100_Valid_Out & channel14_Kernel100_Valid_Out & channel15_Kernel100_Valid_Out & channel16_Kernel100_Valid_Out & channel17_Kernel100_Valid_Out & channel18_Kernel100_Valid_Out & channel19_Kernel100_Valid_Out & channel20_Kernel100_Valid_Out & channel21_Kernel100_Valid_Out & channel22_Kernel100_Valid_Out & channel23_Kernel100_Valid_Out & channel24_Kernel100_Valid_Out & channel25_Kernel100_Valid_Out & channel26_Kernel100_Valid_Out & channel27_Kernel100_Valid_Out & channel28_Kernel100_Valid_Out & channel29_Kernel100_Valid_Out & channel30_Kernel100_Valid_Out & channel31_Kernel100_Valid_Out & channel32_Kernel100_Valid_Out & channel33_Kernel100_Valid_Out & channel34_Kernel100_Valid_Out & channel35_Kernel100_Valid_Out & channel36_Kernel100_Valid_Out & channel37_Kernel100_Valid_Out & channel38_Kernel100_Valid_Out & channel39_Kernel100_Valid_Out & channel40_Kernel100_Valid_Out & channel41_Kernel100_Valid_Out & channel42_Kernel100_Valid_Out & channel43_Kernel100_Valid_Out & channel44_Kernel100_Valid_Out & channel45_Kernel100_Valid_Out & channel46_Kernel100_Valid_Out & channel47_Kernel100_Valid_Out & channel48_Kernel100_Valid_Out & channel49_Kernel100_Valid_Out & channel50_Kernel100_Valid_Out & channel51_Kernel100_Valid_Out & channel52_Kernel100_Valid_Out & channel53_Kernel100_Valid_Out & channel54_Kernel100_Valid_Out & channel55_Kernel100_Valid_Out & channel56_Kernel100_Valid_Out & channel57_Kernel100_Valid_Out & channel58_Kernel100_Valid_Out & channel59_Kernel100_Valid_Out & channel60_Kernel100_Valid_Out & channel61_Kernel100_Valid_Out & channel62_Kernel100_Valid_Out & channel63_Kernel100_Valid_Out & channel64_Kernel100_Valid_Out;

	wire channel1_Kernel101_Valid_Out, channel2_Kernel101_Valid_Out, channel3_Kernel101_Valid_Out, channel4_Kernel101_Valid_Out, channel5_Kernel101_Valid_Out, channel6_Kernel101_Valid_Out, channel7_Kernel101_Valid_Out, channel8_Kernel101_Valid_Out, channel9_Kernel101_Valid_Out, channel10_Kernel101_Valid_Out, channel11_Kernel101_Valid_Out, channel12_Kernel101_Valid_Out, channel13_Kernel101_Valid_Out, channel14_Kernel101_Valid_Out, channel15_Kernel101_Valid_Out, channel16_Kernel101_Valid_Out, channel17_Kernel101_Valid_Out, channel18_Kernel101_Valid_Out, channel19_Kernel101_Valid_Out, channel20_Kernel101_Valid_Out, channel21_Kernel101_Valid_Out, channel22_Kernel101_Valid_Out, channel23_Kernel101_Valid_Out, channel24_Kernel101_Valid_Out, channel25_Kernel101_Valid_Out, channel26_Kernel101_Valid_Out, channel27_Kernel101_Valid_Out, channel28_Kernel101_Valid_Out, channel29_Kernel101_Valid_Out, channel30_Kernel101_Valid_Out, channel31_Kernel101_Valid_Out, channel32_Kernel101_Valid_Out, channel33_Kernel101_Valid_Out, channel34_Kernel101_Valid_Out, channel35_Kernel101_Valid_Out, channel36_Kernel101_Valid_Out, channel37_Kernel101_Valid_Out, channel38_Kernel101_Valid_Out, channel39_Kernel101_Valid_Out, channel40_Kernel101_Valid_Out, channel41_Kernel101_Valid_Out, channel42_Kernel101_Valid_Out, channel43_Kernel101_Valid_Out, channel44_Kernel101_Valid_Out, channel45_Kernel101_Valid_Out, channel46_Kernel101_Valid_Out, channel47_Kernel101_Valid_Out, channel48_Kernel101_Valid_Out, channel49_Kernel101_Valid_Out, channel50_Kernel101_Valid_Out, channel51_Kernel101_Valid_Out, channel52_Kernel101_Valid_Out, channel53_Kernel101_Valid_Out, channel54_Kernel101_Valid_Out, channel55_Kernel101_Valid_Out, channel56_Kernel101_Valid_Out, channel57_Kernel101_Valid_Out, channel58_Kernel101_Valid_Out, channel59_Kernel101_Valid_Out, channel60_Kernel101_Valid_Out, channel61_Kernel101_Valid_Out, channel62_Kernel101_Valid_Out, channel63_Kernel101_Valid_Out, channel64_Kernel101_Valid_Out;

	assign add_kernel101=channel1_Kernel101_Valid_Out & channel2_Kernel101_Valid_Out & channel3_Kernel101_Valid_Out & channel4_Kernel101_Valid_Out & channel5_Kernel101_Valid_Out & channel6_Kernel101_Valid_Out & channel7_Kernel101_Valid_Out & channel8_Kernel101_Valid_Out & channel9_Kernel101_Valid_Out & channel10_Kernel101_Valid_Out & channel11_Kernel101_Valid_Out & channel12_Kernel101_Valid_Out & channel13_Kernel101_Valid_Out & channel14_Kernel101_Valid_Out & channel15_Kernel101_Valid_Out & channel16_Kernel101_Valid_Out & channel17_Kernel101_Valid_Out & channel18_Kernel101_Valid_Out & channel19_Kernel101_Valid_Out & channel20_Kernel101_Valid_Out & channel21_Kernel101_Valid_Out & channel22_Kernel101_Valid_Out & channel23_Kernel101_Valid_Out & channel24_Kernel101_Valid_Out & channel25_Kernel101_Valid_Out & channel26_Kernel101_Valid_Out & channel27_Kernel101_Valid_Out & channel28_Kernel101_Valid_Out & channel29_Kernel101_Valid_Out & channel30_Kernel101_Valid_Out & channel31_Kernel101_Valid_Out & channel32_Kernel101_Valid_Out & channel33_Kernel101_Valid_Out & channel34_Kernel101_Valid_Out & channel35_Kernel101_Valid_Out & channel36_Kernel101_Valid_Out & channel37_Kernel101_Valid_Out & channel38_Kernel101_Valid_Out & channel39_Kernel101_Valid_Out & channel40_Kernel101_Valid_Out & channel41_Kernel101_Valid_Out & channel42_Kernel101_Valid_Out & channel43_Kernel101_Valid_Out & channel44_Kernel101_Valid_Out & channel45_Kernel101_Valid_Out & channel46_Kernel101_Valid_Out & channel47_Kernel101_Valid_Out & channel48_Kernel101_Valid_Out & channel49_Kernel101_Valid_Out & channel50_Kernel101_Valid_Out & channel51_Kernel101_Valid_Out & channel52_Kernel101_Valid_Out & channel53_Kernel101_Valid_Out & channel54_Kernel101_Valid_Out & channel55_Kernel101_Valid_Out & channel56_Kernel101_Valid_Out & channel57_Kernel101_Valid_Out & channel58_Kernel101_Valid_Out & channel59_Kernel101_Valid_Out & channel60_Kernel101_Valid_Out & channel61_Kernel101_Valid_Out & channel62_Kernel101_Valid_Out & channel63_Kernel101_Valid_Out & channel64_Kernel101_Valid_Out;

	wire channel1_Kernel102_Valid_Out, channel2_Kernel102_Valid_Out, channel3_Kernel102_Valid_Out, channel4_Kernel102_Valid_Out, channel5_Kernel102_Valid_Out, channel6_Kernel102_Valid_Out, channel7_Kernel102_Valid_Out, channel8_Kernel102_Valid_Out, channel9_Kernel102_Valid_Out, channel10_Kernel102_Valid_Out, channel11_Kernel102_Valid_Out, channel12_Kernel102_Valid_Out, channel13_Kernel102_Valid_Out, channel14_Kernel102_Valid_Out, channel15_Kernel102_Valid_Out, channel16_Kernel102_Valid_Out, channel17_Kernel102_Valid_Out, channel18_Kernel102_Valid_Out, channel19_Kernel102_Valid_Out, channel20_Kernel102_Valid_Out, channel21_Kernel102_Valid_Out, channel22_Kernel102_Valid_Out, channel23_Kernel102_Valid_Out, channel24_Kernel102_Valid_Out, channel25_Kernel102_Valid_Out, channel26_Kernel102_Valid_Out, channel27_Kernel102_Valid_Out, channel28_Kernel102_Valid_Out, channel29_Kernel102_Valid_Out, channel30_Kernel102_Valid_Out, channel31_Kernel102_Valid_Out, channel32_Kernel102_Valid_Out, channel33_Kernel102_Valid_Out, channel34_Kernel102_Valid_Out, channel35_Kernel102_Valid_Out, channel36_Kernel102_Valid_Out, channel37_Kernel102_Valid_Out, channel38_Kernel102_Valid_Out, channel39_Kernel102_Valid_Out, channel40_Kernel102_Valid_Out, channel41_Kernel102_Valid_Out, channel42_Kernel102_Valid_Out, channel43_Kernel102_Valid_Out, channel44_Kernel102_Valid_Out, channel45_Kernel102_Valid_Out, channel46_Kernel102_Valid_Out, channel47_Kernel102_Valid_Out, channel48_Kernel102_Valid_Out, channel49_Kernel102_Valid_Out, channel50_Kernel102_Valid_Out, channel51_Kernel102_Valid_Out, channel52_Kernel102_Valid_Out, channel53_Kernel102_Valid_Out, channel54_Kernel102_Valid_Out, channel55_Kernel102_Valid_Out, channel56_Kernel102_Valid_Out, channel57_Kernel102_Valid_Out, channel58_Kernel102_Valid_Out, channel59_Kernel102_Valid_Out, channel60_Kernel102_Valid_Out, channel61_Kernel102_Valid_Out, channel62_Kernel102_Valid_Out, channel63_Kernel102_Valid_Out, channel64_Kernel102_Valid_Out;

	assign add_kernel102=channel1_Kernel102_Valid_Out & channel2_Kernel102_Valid_Out & channel3_Kernel102_Valid_Out & channel4_Kernel102_Valid_Out & channel5_Kernel102_Valid_Out & channel6_Kernel102_Valid_Out & channel7_Kernel102_Valid_Out & channel8_Kernel102_Valid_Out & channel9_Kernel102_Valid_Out & channel10_Kernel102_Valid_Out & channel11_Kernel102_Valid_Out & channel12_Kernel102_Valid_Out & channel13_Kernel102_Valid_Out & channel14_Kernel102_Valid_Out & channel15_Kernel102_Valid_Out & channel16_Kernel102_Valid_Out & channel17_Kernel102_Valid_Out & channel18_Kernel102_Valid_Out & channel19_Kernel102_Valid_Out & channel20_Kernel102_Valid_Out & channel21_Kernel102_Valid_Out & channel22_Kernel102_Valid_Out & channel23_Kernel102_Valid_Out & channel24_Kernel102_Valid_Out & channel25_Kernel102_Valid_Out & channel26_Kernel102_Valid_Out & channel27_Kernel102_Valid_Out & channel28_Kernel102_Valid_Out & channel29_Kernel102_Valid_Out & channel30_Kernel102_Valid_Out & channel31_Kernel102_Valid_Out & channel32_Kernel102_Valid_Out & channel33_Kernel102_Valid_Out & channel34_Kernel102_Valid_Out & channel35_Kernel102_Valid_Out & channel36_Kernel102_Valid_Out & channel37_Kernel102_Valid_Out & channel38_Kernel102_Valid_Out & channel39_Kernel102_Valid_Out & channel40_Kernel102_Valid_Out & channel41_Kernel102_Valid_Out & channel42_Kernel102_Valid_Out & channel43_Kernel102_Valid_Out & channel44_Kernel102_Valid_Out & channel45_Kernel102_Valid_Out & channel46_Kernel102_Valid_Out & channel47_Kernel102_Valid_Out & channel48_Kernel102_Valid_Out & channel49_Kernel102_Valid_Out & channel50_Kernel102_Valid_Out & channel51_Kernel102_Valid_Out & channel52_Kernel102_Valid_Out & channel53_Kernel102_Valid_Out & channel54_Kernel102_Valid_Out & channel55_Kernel102_Valid_Out & channel56_Kernel102_Valid_Out & channel57_Kernel102_Valid_Out & channel58_Kernel102_Valid_Out & channel59_Kernel102_Valid_Out & channel60_Kernel102_Valid_Out & channel61_Kernel102_Valid_Out & channel62_Kernel102_Valid_Out & channel63_Kernel102_Valid_Out & channel64_Kernel102_Valid_Out;

	wire channel1_Kernel103_Valid_Out, channel2_Kernel103_Valid_Out, channel3_Kernel103_Valid_Out, channel4_Kernel103_Valid_Out, channel5_Kernel103_Valid_Out, channel6_Kernel103_Valid_Out, channel7_Kernel103_Valid_Out, channel8_Kernel103_Valid_Out, channel9_Kernel103_Valid_Out, channel10_Kernel103_Valid_Out, channel11_Kernel103_Valid_Out, channel12_Kernel103_Valid_Out, channel13_Kernel103_Valid_Out, channel14_Kernel103_Valid_Out, channel15_Kernel103_Valid_Out, channel16_Kernel103_Valid_Out, channel17_Kernel103_Valid_Out, channel18_Kernel103_Valid_Out, channel19_Kernel103_Valid_Out, channel20_Kernel103_Valid_Out, channel21_Kernel103_Valid_Out, channel22_Kernel103_Valid_Out, channel23_Kernel103_Valid_Out, channel24_Kernel103_Valid_Out, channel25_Kernel103_Valid_Out, channel26_Kernel103_Valid_Out, channel27_Kernel103_Valid_Out, channel28_Kernel103_Valid_Out, channel29_Kernel103_Valid_Out, channel30_Kernel103_Valid_Out, channel31_Kernel103_Valid_Out, channel32_Kernel103_Valid_Out, channel33_Kernel103_Valid_Out, channel34_Kernel103_Valid_Out, channel35_Kernel103_Valid_Out, channel36_Kernel103_Valid_Out, channel37_Kernel103_Valid_Out, channel38_Kernel103_Valid_Out, channel39_Kernel103_Valid_Out, channel40_Kernel103_Valid_Out, channel41_Kernel103_Valid_Out, channel42_Kernel103_Valid_Out, channel43_Kernel103_Valid_Out, channel44_Kernel103_Valid_Out, channel45_Kernel103_Valid_Out, channel46_Kernel103_Valid_Out, channel47_Kernel103_Valid_Out, channel48_Kernel103_Valid_Out, channel49_Kernel103_Valid_Out, channel50_Kernel103_Valid_Out, channel51_Kernel103_Valid_Out, channel52_Kernel103_Valid_Out, channel53_Kernel103_Valid_Out, channel54_Kernel103_Valid_Out, channel55_Kernel103_Valid_Out, channel56_Kernel103_Valid_Out, channel57_Kernel103_Valid_Out, channel58_Kernel103_Valid_Out, channel59_Kernel103_Valid_Out, channel60_Kernel103_Valid_Out, channel61_Kernel103_Valid_Out, channel62_Kernel103_Valid_Out, channel63_Kernel103_Valid_Out, channel64_Kernel103_Valid_Out;

	assign add_kernel103=channel1_Kernel103_Valid_Out & channel2_Kernel103_Valid_Out & channel3_Kernel103_Valid_Out & channel4_Kernel103_Valid_Out & channel5_Kernel103_Valid_Out & channel6_Kernel103_Valid_Out & channel7_Kernel103_Valid_Out & channel8_Kernel103_Valid_Out & channel9_Kernel103_Valid_Out & channel10_Kernel103_Valid_Out & channel11_Kernel103_Valid_Out & channel12_Kernel103_Valid_Out & channel13_Kernel103_Valid_Out & channel14_Kernel103_Valid_Out & channel15_Kernel103_Valid_Out & channel16_Kernel103_Valid_Out & channel17_Kernel103_Valid_Out & channel18_Kernel103_Valid_Out & channel19_Kernel103_Valid_Out & channel20_Kernel103_Valid_Out & channel21_Kernel103_Valid_Out & channel22_Kernel103_Valid_Out & channel23_Kernel103_Valid_Out & channel24_Kernel103_Valid_Out & channel25_Kernel103_Valid_Out & channel26_Kernel103_Valid_Out & channel27_Kernel103_Valid_Out & channel28_Kernel103_Valid_Out & channel29_Kernel103_Valid_Out & channel30_Kernel103_Valid_Out & channel31_Kernel103_Valid_Out & channel32_Kernel103_Valid_Out & channel33_Kernel103_Valid_Out & channel34_Kernel103_Valid_Out & channel35_Kernel103_Valid_Out & channel36_Kernel103_Valid_Out & channel37_Kernel103_Valid_Out & channel38_Kernel103_Valid_Out & channel39_Kernel103_Valid_Out & channel40_Kernel103_Valid_Out & channel41_Kernel103_Valid_Out & channel42_Kernel103_Valid_Out & channel43_Kernel103_Valid_Out & channel44_Kernel103_Valid_Out & channel45_Kernel103_Valid_Out & channel46_Kernel103_Valid_Out & channel47_Kernel103_Valid_Out & channel48_Kernel103_Valid_Out & channel49_Kernel103_Valid_Out & channel50_Kernel103_Valid_Out & channel51_Kernel103_Valid_Out & channel52_Kernel103_Valid_Out & channel53_Kernel103_Valid_Out & channel54_Kernel103_Valid_Out & channel55_Kernel103_Valid_Out & channel56_Kernel103_Valid_Out & channel57_Kernel103_Valid_Out & channel58_Kernel103_Valid_Out & channel59_Kernel103_Valid_Out & channel60_Kernel103_Valid_Out & channel61_Kernel103_Valid_Out & channel62_Kernel103_Valid_Out & channel63_Kernel103_Valid_Out & channel64_Kernel103_Valid_Out;

	wire channel1_Kernel104_Valid_Out, channel2_Kernel104_Valid_Out, channel3_Kernel104_Valid_Out, channel4_Kernel104_Valid_Out, channel5_Kernel104_Valid_Out, channel6_Kernel104_Valid_Out, channel7_Kernel104_Valid_Out, channel8_Kernel104_Valid_Out, channel9_Kernel104_Valid_Out, channel10_Kernel104_Valid_Out, channel11_Kernel104_Valid_Out, channel12_Kernel104_Valid_Out, channel13_Kernel104_Valid_Out, channel14_Kernel104_Valid_Out, channel15_Kernel104_Valid_Out, channel16_Kernel104_Valid_Out, channel17_Kernel104_Valid_Out, channel18_Kernel104_Valid_Out, channel19_Kernel104_Valid_Out, channel20_Kernel104_Valid_Out, channel21_Kernel104_Valid_Out, channel22_Kernel104_Valid_Out, channel23_Kernel104_Valid_Out, channel24_Kernel104_Valid_Out, channel25_Kernel104_Valid_Out, channel26_Kernel104_Valid_Out, channel27_Kernel104_Valid_Out, channel28_Kernel104_Valid_Out, channel29_Kernel104_Valid_Out, channel30_Kernel104_Valid_Out, channel31_Kernel104_Valid_Out, channel32_Kernel104_Valid_Out, channel33_Kernel104_Valid_Out, channel34_Kernel104_Valid_Out, channel35_Kernel104_Valid_Out, channel36_Kernel104_Valid_Out, channel37_Kernel104_Valid_Out, channel38_Kernel104_Valid_Out, channel39_Kernel104_Valid_Out, channel40_Kernel104_Valid_Out, channel41_Kernel104_Valid_Out, channel42_Kernel104_Valid_Out, channel43_Kernel104_Valid_Out, channel44_Kernel104_Valid_Out, channel45_Kernel104_Valid_Out, channel46_Kernel104_Valid_Out, channel47_Kernel104_Valid_Out, channel48_Kernel104_Valid_Out, channel49_Kernel104_Valid_Out, channel50_Kernel104_Valid_Out, channel51_Kernel104_Valid_Out, channel52_Kernel104_Valid_Out, channel53_Kernel104_Valid_Out, channel54_Kernel104_Valid_Out, channel55_Kernel104_Valid_Out, channel56_Kernel104_Valid_Out, channel57_Kernel104_Valid_Out, channel58_Kernel104_Valid_Out, channel59_Kernel104_Valid_Out, channel60_Kernel104_Valid_Out, channel61_Kernel104_Valid_Out, channel62_Kernel104_Valid_Out, channel63_Kernel104_Valid_Out, channel64_Kernel104_Valid_Out;

	assign add_kernel104=channel1_Kernel104_Valid_Out & channel2_Kernel104_Valid_Out & channel3_Kernel104_Valid_Out & channel4_Kernel104_Valid_Out & channel5_Kernel104_Valid_Out & channel6_Kernel104_Valid_Out & channel7_Kernel104_Valid_Out & channel8_Kernel104_Valid_Out & channel9_Kernel104_Valid_Out & channel10_Kernel104_Valid_Out & channel11_Kernel104_Valid_Out & channel12_Kernel104_Valid_Out & channel13_Kernel104_Valid_Out & channel14_Kernel104_Valid_Out & channel15_Kernel104_Valid_Out & channel16_Kernel104_Valid_Out & channel17_Kernel104_Valid_Out & channel18_Kernel104_Valid_Out & channel19_Kernel104_Valid_Out & channel20_Kernel104_Valid_Out & channel21_Kernel104_Valid_Out & channel22_Kernel104_Valid_Out & channel23_Kernel104_Valid_Out & channel24_Kernel104_Valid_Out & channel25_Kernel104_Valid_Out & channel26_Kernel104_Valid_Out & channel27_Kernel104_Valid_Out & channel28_Kernel104_Valid_Out & channel29_Kernel104_Valid_Out & channel30_Kernel104_Valid_Out & channel31_Kernel104_Valid_Out & channel32_Kernel104_Valid_Out & channel33_Kernel104_Valid_Out & channel34_Kernel104_Valid_Out & channel35_Kernel104_Valid_Out & channel36_Kernel104_Valid_Out & channel37_Kernel104_Valid_Out & channel38_Kernel104_Valid_Out & channel39_Kernel104_Valid_Out & channel40_Kernel104_Valid_Out & channel41_Kernel104_Valid_Out & channel42_Kernel104_Valid_Out & channel43_Kernel104_Valid_Out & channel44_Kernel104_Valid_Out & channel45_Kernel104_Valid_Out & channel46_Kernel104_Valid_Out & channel47_Kernel104_Valid_Out & channel48_Kernel104_Valid_Out & channel49_Kernel104_Valid_Out & channel50_Kernel104_Valid_Out & channel51_Kernel104_Valid_Out & channel52_Kernel104_Valid_Out & channel53_Kernel104_Valid_Out & channel54_Kernel104_Valid_Out & channel55_Kernel104_Valid_Out & channel56_Kernel104_Valid_Out & channel57_Kernel104_Valid_Out & channel58_Kernel104_Valid_Out & channel59_Kernel104_Valid_Out & channel60_Kernel104_Valid_Out & channel61_Kernel104_Valid_Out & channel62_Kernel104_Valid_Out & channel63_Kernel104_Valid_Out & channel64_Kernel104_Valid_Out;

	wire channel1_Kernel105_Valid_Out, channel2_Kernel105_Valid_Out, channel3_Kernel105_Valid_Out, channel4_Kernel105_Valid_Out, channel5_Kernel105_Valid_Out, channel6_Kernel105_Valid_Out, channel7_Kernel105_Valid_Out, channel8_Kernel105_Valid_Out, channel9_Kernel105_Valid_Out, channel10_Kernel105_Valid_Out, channel11_Kernel105_Valid_Out, channel12_Kernel105_Valid_Out, channel13_Kernel105_Valid_Out, channel14_Kernel105_Valid_Out, channel15_Kernel105_Valid_Out, channel16_Kernel105_Valid_Out, channel17_Kernel105_Valid_Out, channel18_Kernel105_Valid_Out, channel19_Kernel105_Valid_Out, channel20_Kernel105_Valid_Out, channel21_Kernel105_Valid_Out, channel22_Kernel105_Valid_Out, channel23_Kernel105_Valid_Out, channel24_Kernel105_Valid_Out, channel25_Kernel105_Valid_Out, channel26_Kernel105_Valid_Out, channel27_Kernel105_Valid_Out, channel28_Kernel105_Valid_Out, channel29_Kernel105_Valid_Out, channel30_Kernel105_Valid_Out, channel31_Kernel105_Valid_Out, channel32_Kernel105_Valid_Out, channel33_Kernel105_Valid_Out, channel34_Kernel105_Valid_Out, channel35_Kernel105_Valid_Out, channel36_Kernel105_Valid_Out, channel37_Kernel105_Valid_Out, channel38_Kernel105_Valid_Out, channel39_Kernel105_Valid_Out, channel40_Kernel105_Valid_Out, channel41_Kernel105_Valid_Out, channel42_Kernel105_Valid_Out, channel43_Kernel105_Valid_Out, channel44_Kernel105_Valid_Out, channel45_Kernel105_Valid_Out, channel46_Kernel105_Valid_Out, channel47_Kernel105_Valid_Out, channel48_Kernel105_Valid_Out, channel49_Kernel105_Valid_Out, channel50_Kernel105_Valid_Out, channel51_Kernel105_Valid_Out, channel52_Kernel105_Valid_Out, channel53_Kernel105_Valid_Out, channel54_Kernel105_Valid_Out, channel55_Kernel105_Valid_Out, channel56_Kernel105_Valid_Out, channel57_Kernel105_Valid_Out, channel58_Kernel105_Valid_Out, channel59_Kernel105_Valid_Out, channel60_Kernel105_Valid_Out, channel61_Kernel105_Valid_Out, channel62_Kernel105_Valid_Out, channel63_Kernel105_Valid_Out, channel64_Kernel105_Valid_Out;

	assign add_kernel105=channel1_Kernel105_Valid_Out & channel2_Kernel105_Valid_Out & channel3_Kernel105_Valid_Out & channel4_Kernel105_Valid_Out & channel5_Kernel105_Valid_Out & channel6_Kernel105_Valid_Out & channel7_Kernel105_Valid_Out & channel8_Kernel105_Valid_Out & channel9_Kernel105_Valid_Out & channel10_Kernel105_Valid_Out & channel11_Kernel105_Valid_Out & channel12_Kernel105_Valid_Out & channel13_Kernel105_Valid_Out & channel14_Kernel105_Valid_Out & channel15_Kernel105_Valid_Out & channel16_Kernel105_Valid_Out & channel17_Kernel105_Valid_Out & channel18_Kernel105_Valid_Out & channel19_Kernel105_Valid_Out & channel20_Kernel105_Valid_Out & channel21_Kernel105_Valid_Out & channel22_Kernel105_Valid_Out & channel23_Kernel105_Valid_Out & channel24_Kernel105_Valid_Out & channel25_Kernel105_Valid_Out & channel26_Kernel105_Valid_Out & channel27_Kernel105_Valid_Out & channel28_Kernel105_Valid_Out & channel29_Kernel105_Valid_Out & channel30_Kernel105_Valid_Out & channel31_Kernel105_Valid_Out & channel32_Kernel105_Valid_Out & channel33_Kernel105_Valid_Out & channel34_Kernel105_Valid_Out & channel35_Kernel105_Valid_Out & channel36_Kernel105_Valid_Out & channel37_Kernel105_Valid_Out & channel38_Kernel105_Valid_Out & channel39_Kernel105_Valid_Out & channel40_Kernel105_Valid_Out & channel41_Kernel105_Valid_Out & channel42_Kernel105_Valid_Out & channel43_Kernel105_Valid_Out & channel44_Kernel105_Valid_Out & channel45_Kernel105_Valid_Out & channel46_Kernel105_Valid_Out & channel47_Kernel105_Valid_Out & channel48_Kernel105_Valid_Out & channel49_Kernel105_Valid_Out & channel50_Kernel105_Valid_Out & channel51_Kernel105_Valid_Out & channel52_Kernel105_Valid_Out & channel53_Kernel105_Valid_Out & channel54_Kernel105_Valid_Out & channel55_Kernel105_Valid_Out & channel56_Kernel105_Valid_Out & channel57_Kernel105_Valid_Out & channel58_Kernel105_Valid_Out & channel59_Kernel105_Valid_Out & channel60_Kernel105_Valid_Out & channel61_Kernel105_Valid_Out & channel62_Kernel105_Valid_Out & channel63_Kernel105_Valid_Out & channel64_Kernel105_Valid_Out;

	wire channel1_Kernel106_Valid_Out, channel2_Kernel106_Valid_Out, channel3_Kernel106_Valid_Out, channel4_Kernel106_Valid_Out, channel5_Kernel106_Valid_Out, channel6_Kernel106_Valid_Out, channel7_Kernel106_Valid_Out, channel8_Kernel106_Valid_Out, channel9_Kernel106_Valid_Out, channel10_Kernel106_Valid_Out, channel11_Kernel106_Valid_Out, channel12_Kernel106_Valid_Out, channel13_Kernel106_Valid_Out, channel14_Kernel106_Valid_Out, channel15_Kernel106_Valid_Out, channel16_Kernel106_Valid_Out, channel17_Kernel106_Valid_Out, channel18_Kernel106_Valid_Out, channel19_Kernel106_Valid_Out, channel20_Kernel106_Valid_Out, channel21_Kernel106_Valid_Out, channel22_Kernel106_Valid_Out, channel23_Kernel106_Valid_Out, channel24_Kernel106_Valid_Out, channel25_Kernel106_Valid_Out, channel26_Kernel106_Valid_Out, channel27_Kernel106_Valid_Out, channel28_Kernel106_Valid_Out, channel29_Kernel106_Valid_Out, channel30_Kernel106_Valid_Out, channel31_Kernel106_Valid_Out, channel32_Kernel106_Valid_Out, channel33_Kernel106_Valid_Out, channel34_Kernel106_Valid_Out, channel35_Kernel106_Valid_Out, channel36_Kernel106_Valid_Out, channel37_Kernel106_Valid_Out, channel38_Kernel106_Valid_Out, channel39_Kernel106_Valid_Out, channel40_Kernel106_Valid_Out, channel41_Kernel106_Valid_Out, channel42_Kernel106_Valid_Out, channel43_Kernel106_Valid_Out, channel44_Kernel106_Valid_Out, channel45_Kernel106_Valid_Out, channel46_Kernel106_Valid_Out, channel47_Kernel106_Valid_Out, channel48_Kernel106_Valid_Out, channel49_Kernel106_Valid_Out, channel50_Kernel106_Valid_Out, channel51_Kernel106_Valid_Out, channel52_Kernel106_Valid_Out, channel53_Kernel106_Valid_Out, channel54_Kernel106_Valid_Out, channel55_Kernel106_Valid_Out, channel56_Kernel106_Valid_Out, channel57_Kernel106_Valid_Out, channel58_Kernel106_Valid_Out, channel59_Kernel106_Valid_Out, channel60_Kernel106_Valid_Out, channel61_Kernel106_Valid_Out, channel62_Kernel106_Valid_Out, channel63_Kernel106_Valid_Out, channel64_Kernel106_Valid_Out;

	assign add_kernel106=channel1_Kernel106_Valid_Out & channel2_Kernel106_Valid_Out & channel3_Kernel106_Valid_Out & channel4_Kernel106_Valid_Out & channel5_Kernel106_Valid_Out & channel6_Kernel106_Valid_Out & channel7_Kernel106_Valid_Out & channel8_Kernel106_Valid_Out & channel9_Kernel106_Valid_Out & channel10_Kernel106_Valid_Out & channel11_Kernel106_Valid_Out & channel12_Kernel106_Valid_Out & channel13_Kernel106_Valid_Out & channel14_Kernel106_Valid_Out & channel15_Kernel106_Valid_Out & channel16_Kernel106_Valid_Out & channel17_Kernel106_Valid_Out & channel18_Kernel106_Valid_Out & channel19_Kernel106_Valid_Out & channel20_Kernel106_Valid_Out & channel21_Kernel106_Valid_Out & channel22_Kernel106_Valid_Out & channel23_Kernel106_Valid_Out & channel24_Kernel106_Valid_Out & channel25_Kernel106_Valid_Out & channel26_Kernel106_Valid_Out & channel27_Kernel106_Valid_Out & channel28_Kernel106_Valid_Out & channel29_Kernel106_Valid_Out & channel30_Kernel106_Valid_Out & channel31_Kernel106_Valid_Out & channel32_Kernel106_Valid_Out & channel33_Kernel106_Valid_Out & channel34_Kernel106_Valid_Out & channel35_Kernel106_Valid_Out & channel36_Kernel106_Valid_Out & channel37_Kernel106_Valid_Out & channel38_Kernel106_Valid_Out & channel39_Kernel106_Valid_Out & channel40_Kernel106_Valid_Out & channel41_Kernel106_Valid_Out & channel42_Kernel106_Valid_Out & channel43_Kernel106_Valid_Out & channel44_Kernel106_Valid_Out & channel45_Kernel106_Valid_Out & channel46_Kernel106_Valid_Out & channel47_Kernel106_Valid_Out & channel48_Kernel106_Valid_Out & channel49_Kernel106_Valid_Out & channel50_Kernel106_Valid_Out & channel51_Kernel106_Valid_Out & channel52_Kernel106_Valid_Out & channel53_Kernel106_Valid_Out & channel54_Kernel106_Valid_Out & channel55_Kernel106_Valid_Out & channel56_Kernel106_Valid_Out & channel57_Kernel106_Valid_Out & channel58_Kernel106_Valid_Out & channel59_Kernel106_Valid_Out & channel60_Kernel106_Valid_Out & channel61_Kernel106_Valid_Out & channel62_Kernel106_Valid_Out & channel63_Kernel106_Valid_Out & channel64_Kernel106_Valid_Out;

	wire channel1_Kernel107_Valid_Out, channel2_Kernel107_Valid_Out, channel3_Kernel107_Valid_Out, channel4_Kernel107_Valid_Out, channel5_Kernel107_Valid_Out, channel6_Kernel107_Valid_Out, channel7_Kernel107_Valid_Out, channel8_Kernel107_Valid_Out, channel9_Kernel107_Valid_Out, channel10_Kernel107_Valid_Out, channel11_Kernel107_Valid_Out, channel12_Kernel107_Valid_Out, channel13_Kernel107_Valid_Out, channel14_Kernel107_Valid_Out, channel15_Kernel107_Valid_Out, channel16_Kernel107_Valid_Out, channel17_Kernel107_Valid_Out, channel18_Kernel107_Valid_Out, channel19_Kernel107_Valid_Out, channel20_Kernel107_Valid_Out, channel21_Kernel107_Valid_Out, channel22_Kernel107_Valid_Out, channel23_Kernel107_Valid_Out, channel24_Kernel107_Valid_Out, channel25_Kernel107_Valid_Out, channel26_Kernel107_Valid_Out, channel27_Kernel107_Valid_Out, channel28_Kernel107_Valid_Out, channel29_Kernel107_Valid_Out, channel30_Kernel107_Valid_Out, channel31_Kernel107_Valid_Out, channel32_Kernel107_Valid_Out, channel33_Kernel107_Valid_Out, channel34_Kernel107_Valid_Out, channel35_Kernel107_Valid_Out, channel36_Kernel107_Valid_Out, channel37_Kernel107_Valid_Out, channel38_Kernel107_Valid_Out, channel39_Kernel107_Valid_Out, channel40_Kernel107_Valid_Out, channel41_Kernel107_Valid_Out, channel42_Kernel107_Valid_Out, channel43_Kernel107_Valid_Out, channel44_Kernel107_Valid_Out, channel45_Kernel107_Valid_Out, channel46_Kernel107_Valid_Out, channel47_Kernel107_Valid_Out, channel48_Kernel107_Valid_Out, channel49_Kernel107_Valid_Out, channel50_Kernel107_Valid_Out, channel51_Kernel107_Valid_Out, channel52_Kernel107_Valid_Out, channel53_Kernel107_Valid_Out, channel54_Kernel107_Valid_Out, channel55_Kernel107_Valid_Out, channel56_Kernel107_Valid_Out, channel57_Kernel107_Valid_Out, channel58_Kernel107_Valid_Out, channel59_Kernel107_Valid_Out, channel60_Kernel107_Valid_Out, channel61_Kernel107_Valid_Out, channel62_Kernel107_Valid_Out, channel63_Kernel107_Valid_Out, channel64_Kernel107_Valid_Out;

	assign add_kernel107=channel1_Kernel107_Valid_Out & channel2_Kernel107_Valid_Out & channel3_Kernel107_Valid_Out & channel4_Kernel107_Valid_Out & channel5_Kernel107_Valid_Out & channel6_Kernel107_Valid_Out & channel7_Kernel107_Valid_Out & channel8_Kernel107_Valid_Out & channel9_Kernel107_Valid_Out & channel10_Kernel107_Valid_Out & channel11_Kernel107_Valid_Out & channel12_Kernel107_Valid_Out & channel13_Kernel107_Valid_Out & channel14_Kernel107_Valid_Out & channel15_Kernel107_Valid_Out & channel16_Kernel107_Valid_Out & channel17_Kernel107_Valid_Out & channel18_Kernel107_Valid_Out & channel19_Kernel107_Valid_Out & channel20_Kernel107_Valid_Out & channel21_Kernel107_Valid_Out & channel22_Kernel107_Valid_Out & channel23_Kernel107_Valid_Out & channel24_Kernel107_Valid_Out & channel25_Kernel107_Valid_Out & channel26_Kernel107_Valid_Out & channel27_Kernel107_Valid_Out & channel28_Kernel107_Valid_Out & channel29_Kernel107_Valid_Out & channel30_Kernel107_Valid_Out & channel31_Kernel107_Valid_Out & channel32_Kernel107_Valid_Out & channel33_Kernel107_Valid_Out & channel34_Kernel107_Valid_Out & channel35_Kernel107_Valid_Out & channel36_Kernel107_Valid_Out & channel37_Kernel107_Valid_Out & channel38_Kernel107_Valid_Out & channel39_Kernel107_Valid_Out & channel40_Kernel107_Valid_Out & channel41_Kernel107_Valid_Out & channel42_Kernel107_Valid_Out & channel43_Kernel107_Valid_Out & channel44_Kernel107_Valid_Out & channel45_Kernel107_Valid_Out & channel46_Kernel107_Valid_Out & channel47_Kernel107_Valid_Out & channel48_Kernel107_Valid_Out & channel49_Kernel107_Valid_Out & channel50_Kernel107_Valid_Out & channel51_Kernel107_Valid_Out & channel52_Kernel107_Valid_Out & channel53_Kernel107_Valid_Out & channel54_Kernel107_Valid_Out & channel55_Kernel107_Valid_Out & channel56_Kernel107_Valid_Out & channel57_Kernel107_Valid_Out & channel58_Kernel107_Valid_Out & channel59_Kernel107_Valid_Out & channel60_Kernel107_Valid_Out & channel61_Kernel107_Valid_Out & channel62_Kernel107_Valid_Out & channel63_Kernel107_Valid_Out & channel64_Kernel107_Valid_Out;

	wire channel1_Kernel108_Valid_Out, channel2_Kernel108_Valid_Out, channel3_Kernel108_Valid_Out, channel4_Kernel108_Valid_Out, channel5_Kernel108_Valid_Out, channel6_Kernel108_Valid_Out, channel7_Kernel108_Valid_Out, channel8_Kernel108_Valid_Out, channel9_Kernel108_Valid_Out, channel10_Kernel108_Valid_Out, channel11_Kernel108_Valid_Out, channel12_Kernel108_Valid_Out, channel13_Kernel108_Valid_Out, channel14_Kernel108_Valid_Out, channel15_Kernel108_Valid_Out, channel16_Kernel108_Valid_Out, channel17_Kernel108_Valid_Out, channel18_Kernel108_Valid_Out, channel19_Kernel108_Valid_Out, channel20_Kernel108_Valid_Out, channel21_Kernel108_Valid_Out, channel22_Kernel108_Valid_Out, channel23_Kernel108_Valid_Out, channel24_Kernel108_Valid_Out, channel25_Kernel108_Valid_Out, channel26_Kernel108_Valid_Out, channel27_Kernel108_Valid_Out, channel28_Kernel108_Valid_Out, channel29_Kernel108_Valid_Out, channel30_Kernel108_Valid_Out, channel31_Kernel108_Valid_Out, channel32_Kernel108_Valid_Out, channel33_Kernel108_Valid_Out, channel34_Kernel108_Valid_Out, channel35_Kernel108_Valid_Out, channel36_Kernel108_Valid_Out, channel37_Kernel108_Valid_Out, channel38_Kernel108_Valid_Out, channel39_Kernel108_Valid_Out, channel40_Kernel108_Valid_Out, channel41_Kernel108_Valid_Out, channel42_Kernel108_Valid_Out, channel43_Kernel108_Valid_Out, channel44_Kernel108_Valid_Out, channel45_Kernel108_Valid_Out, channel46_Kernel108_Valid_Out, channel47_Kernel108_Valid_Out, channel48_Kernel108_Valid_Out, channel49_Kernel108_Valid_Out, channel50_Kernel108_Valid_Out, channel51_Kernel108_Valid_Out, channel52_Kernel108_Valid_Out, channel53_Kernel108_Valid_Out, channel54_Kernel108_Valid_Out, channel55_Kernel108_Valid_Out, channel56_Kernel108_Valid_Out, channel57_Kernel108_Valid_Out, channel58_Kernel108_Valid_Out, channel59_Kernel108_Valid_Out, channel60_Kernel108_Valid_Out, channel61_Kernel108_Valid_Out, channel62_Kernel108_Valid_Out, channel63_Kernel108_Valid_Out, channel64_Kernel108_Valid_Out;

	assign add_kernel108=channel1_Kernel108_Valid_Out & channel2_Kernel108_Valid_Out & channel3_Kernel108_Valid_Out & channel4_Kernel108_Valid_Out & channel5_Kernel108_Valid_Out & channel6_Kernel108_Valid_Out & channel7_Kernel108_Valid_Out & channel8_Kernel108_Valid_Out & channel9_Kernel108_Valid_Out & channel10_Kernel108_Valid_Out & channel11_Kernel108_Valid_Out & channel12_Kernel108_Valid_Out & channel13_Kernel108_Valid_Out & channel14_Kernel108_Valid_Out & channel15_Kernel108_Valid_Out & channel16_Kernel108_Valid_Out & channel17_Kernel108_Valid_Out & channel18_Kernel108_Valid_Out & channel19_Kernel108_Valid_Out & channel20_Kernel108_Valid_Out & channel21_Kernel108_Valid_Out & channel22_Kernel108_Valid_Out & channel23_Kernel108_Valid_Out & channel24_Kernel108_Valid_Out & channel25_Kernel108_Valid_Out & channel26_Kernel108_Valid_Out & channel27_Kernel108_Valid_Out & channel28_Kernel108_Valid_Out & channel29_Kernel108_Valid_Out & channel30_Kernel108_Valid_Out & channel31_Kernel108_Valid_Out & channel32_Kernel108_Valid_Out & channel33_Kernel108_Valid_Out & channel34_Kernel108_Valid_Out & channel35_Kernel108_Valid_Out & channel36_Kernel108_Valid_Out & channel37_Kernel108_Valid_Out & channel38_Kernel108_Valid_Out & channel39_Kernel108_Valid_Out & channel40_Kernel108_Valid_Out & channel41_Kernel108_Valid_Out & channel42_Kernel108_Valid_Out & channel43_Kernel108_Valid_Out & channel44_Kernel108_Valid_Out & channel45_Kernel108_Valid_Out & channel46_Kernel108_Valid_Out & channel47_Kernel108_Valid_Out & channel48_Kernel108_Valid_Out & channel49_Kernel108_Valid_Out & channel50_Kernel108_Valid_Out & channel51_Kernel108_Valid_Out & channel52_Kernel108_Valid_Out & channel53_Kernel108_Valid_Out & channel54_Kernel108_Valid_Out & channel55_Kernel108_Valid_Out & channel56_Kernel108_Valid_Out & channel57_Kernel108_Valid_Out & channel58_Kernel108_Valid_Out & channel59_Kernel108_Valid_Out & channel60_Kernel108_Valid_Out & channel61_Kernel108_Valid_Out & channel62_Kernel108_Valid_Out & channel63_Kernel108_Valid_Out & channel64_Kernel108_Valid_Out;

	wire channel1_Kernel109_Valid_Out, channel2_Kernel109_Valid_Out, channel3_Kernel109_Valid_Out, channel4_Kernel109_Valid_Out, channel5_Kernel109_Valid_Out, channel6_Kernel109_Valid_Out, channel7_Kernel109_Valid_Out, channel8_Kernel109_Valid_Out, channel9_Kernel109_Valid_Out, channel10_Kernel109_Valid_Out, channel11_Kernel109_Valid_Out, channel12_Kernel109_Valid_Out, channel13_Kernel109_Valid_Out, channel14_Kernel109_Valid_Out, channel15_Kernel109_Valid_Out, channel16_Kernel109_Valid_Out, channel17_Kernel109_Valid_Out, channel18_Kernel109_Valid_Out, channel19_Kernel109_Valid_Out, channel20_Kernel109_Valid_Out, channel21_Kernel109_Valid_Out, channel22_Kernel109_Valid_Out, channel23_Kernel109_Valid_Out, channel24_Kernel109_Valid_Out, channel25_Kernel109_Valid_Out, channel26_Kernel109_Valid_Out, channel27_Kernel109_Valid_Out, channel28_Kernel109_Valid_Out, channel29_Kernel109_Valid_Out, channel30_Kernel109_Valid_Out, channel31_Kernel109_Valid_Out, channel32_Kernel109_Valid_Out, channel33_Kernel109_Valid_Out, channel34_Kernel109_Valid_Out, channel35_Kernel109_Valid_Out, channel36_Kernel109_Valid_Out, channel37_Kernel109_Valid_Out, channel38_Kernel109_Valid_Out, channel39_Kernel109_Valid_Out, channel40_Kernel109_Valid_Out, channel41_Kernel109_Valid_Out, channel42_Kernel109_Valid_Out, channel43_Kernel109_Valid_Out, channel44_Kernel109_Valid_Out, channel45_Kernel109_Valid_Out, channel46_Kernel109_Valid_Out, channel47_Kernel109_Valid_Out, channel48_Kernel109_Valid_Out, channel49_Kernel109_Valid_Out, channel50_Kernel109_Valid_Out, channel51_Kernel109_Valid_Out, channel52_Kernel109_Valid_Out, channel53_Kernel109_Valid_Out, channel54_Kernel109_Valid_Out, channel55_Kernel109_Valid_Out, channel56_Kernel109_Valid_Out, channel57_Kernel109_Valid_Out, channel58_Kernel109_Valid_Out, channel59_Kernel109_Valid_Out, channel60_Kernel109_Valid_Out, channel61_Kernel109_Valid_Out, channel62_Kernel109_Valid_Out, channel63_Kernel109_Valid_Out, channel64_Kernel109_Valid_Out;

	assign add_kernel109=channel1_Kernel109_Valid_Out & channel2_Kernel109_Valid_Out & channel3_Kernel109_Valid_Out & channel4_Kernel109_Valid_Out & channel5_Kernel109_Valid_Out & channel6_Kernel109_Valid_Out & channel7_Kernel109_Valid_Out & channel8_Kernel109_Valid_Out & channel9_Kernel109_Valid_Out & channel10_Kernel109_Valid_Out & channel11_Kernel109_Valid_Out & channel12_Kernel109_Valid_Out & channel13_Kernel109_Valid_Out & channel14_Kernel109_Valid_Out & channel15_Kernel109_Valid_Out & channel16_Kernel109_Valid_Out & channel17_Kernel109_Valid_Out & channel18_Kernel109_Valid_Out & channel19_Kernel109_Valid_Out & channel20_Kernel109_Valid_Out & channel21_Kernel109_Valid_Out & channel22_Kernel109_Valid_Out & channel23_Kernel109_Valid_Out & channel24_Kernel109_Valid_Out & channel25_Kernel109_Valid_Out & channel26_Kernel109_Valid_Out & channel27_Kernel109_Valid_Out & channel28_Kernel109_Valid_Out & channel29_Kernel109_Valid_Out & channel30_Kernel109_Valid_Out & channel31_Kernel109_Valid_Out & channel32_Kernel109_Valid_Out & channel33_Kernel109_Valid_Out & channel34_Kernel109_Valid_Out & channel35_Kernel109_Valid_Out & channel36_Kernel109_Valid_Out & channel37_Kernel109_Valid_Out & channel38_Kernel109_Valid_Out & channel39_Kernel109_Valid_Out & channel40_Kernel109_Valid_Out & channel41_Kernel109_Valid_Out & channel42_Kernel109_Valid_Out & channel43_Kernel109_Valid_Out & channel44_Kernel109_Valid_Out & channel45_Kernel109_Valid_Out & channel46_Kernel109_Valid_Out & channel47_Kernel109_Valid_Out & channel48_Kernel109_Valid_Out & channel49_Kernel109_Valid_Out & channel50_Kernel109_Valid_Out & channel51_Kernel109_Valid_Out & channel52_Kernel109_Valid_Out & channel53_Kernel109_Valid_Out & channel54_Kernel109_Valid_Out & channel55_Kernel109_Valid_Out & channel56_Kernel109_Valid_Out & channel57_Kernel109_Valid_Out & channel58_Kernel109_Valid_Out & channel59_Kernel109_Valid_Out & channel60_Kernel109_Valid_Out & channel61_Kernel109_Valid_Out & channel62_Kernel109_Valid_Out & channel63_Kernel109_Valid_Out & channel64_Kernel109_Valid_Out;

	wire channel1_Kernel110_Valid_Out, channel2_Kernel110_Valid_Out, channel3_Kernel110_Valid_Out, channel4_Kernel110_Valid_Out, channel5_Kernel110_Valid_Out, channel6_Kernel110_Valid_Out, channel7_Kernel110_Valid_Out, channel8_Kernel110_Valid_Out, channel9_Kernel110_Valid_Out, channel10_Kernel110_Valid_Out, channel11_Kernel110_Valid_Out, channel12_Kernel110_Valid_Out, channel13_Kernel110_Valid_Out, channel14_Kernel110_Valid_Out, channel15_Kernel110_Valid_Out, channel16_Kernel110_Valid_Out, channel17_Kernel110_Valid_Out, channel18_Kernel110_Valid_Out, channel19_Kernel110_Valid_Out, channel20_Kernel110_Valid_Out, channel21_Kernel110_Valid_Out, channel22_Kernel110_Valid_Out, channel23_Kernel110_Valid_Out, channel24_Kernel110_Valid_Out, channel25_Kernel110_Valid_Out, channel26_Kernel110_Valid_Out, channel27_Kernel110_Valid_Out, channel28_Kernel110_Valid_Out, channel29_Kernel110_Valid_Out, channel30_Kernel110_Valid_Out, channel31_Kernel110_Valid_Out, channel32_Kernel110_Valid_Out, channel33_Kernel110_Valid_Out, channel34_Kernel110_Valid_Out, channel35_Kernel110_Valid_Out, channel36_Kernel110_Valid_Out, channel37_Kernel110_Valid_Out, channel38_Kernel110_Valid_Out, channel39_Kernel110_Valid_Out, channel40_Kernel110_Valid_Out, channel41_Kernel110_Valid_Out, channel42_Kernel110_Valid_Out, channel43_Kernel110_Valid_Out, channel44_Kernel110_Valid_Out, channel45_Kernel110_Valid_Out, channel46_Kernel110_Valid_Out, channel47_Kernel110_Valid_Out, channel48_Kernel110_Valid_Out, channel49_Kernel110_Valid_Out, channel50_Kernel110_Valid_Out, channel51_Kernel110_Valid_Out, channel52_Kernel110_Valid_Out, channel53_Kernel110_Valid_Out, channel54_Kernel110_Valid_Out, channel55_Kernel110_Valid_Out, channel56_Kernel110_Valid_Out, channel57_Kernel110_Valid_Out, channel58_Kernel110_Valid_Out, channel59_Kernel110_Valid_Out, channel60_Kernel110_Valid_Out, channel61_Kernel110_Valid_Out, channel62_Kernel110_Valid_Out, channel63_Kernel110_Valid_Out, channel64_Kernel110_Valid_Out;

	assign add_kernel110=channel1_Kernel110_Valid_Out & channel2_Kernel110_Valid_Out & channel3_Kernel110_Valid_Out & channel4_Kernel110_Valid_Out & channel5_Kernel110_Valid_Out & channel6_Kernel110_Valid_Out & channel7_Kernel110_Valid_Out & channel8_Kernel110_Valid_Out & channel9_Kernel110_Valid_Out & channel10_Kernel110_Valid_Out & channel11_Kernel110_Valid_Out & channel12_Kernel110_Valid_Out & channel13_Kernel110_Valid_Out & channel14_Kernel110_Valid_Out & channel15_Kernel110_Valid_Out & channel16_Kernel110_Valid_Out & channel17_Kernel110_Valid_Out & channel18_Kernel110_Valid_Out & channel19_Kernel110_Valid_Out & channel20_Kernel110_Valid_Out & channel21_Kernel110_Valid_Out & channel22_Kernel110_Valid_Out & channel23_Kernel110_Valid_Out & channel24_Kernel110_Valid_Out & channel25_Kernel110_Valid_Out & channel26_Kernel110_Valid_Out & channel27_Kernel110_Valid_Out & channel28_Kernel110_Valid_Out & channel29_Kernel110_Valid_Out & channel30_Kernel110_Valid_Out & channel31_Kernel110_Valid_Out & channel32_Kernel110_Valid_Out & channel33_Kernel110_Valid_Out & channel34_Kernel110_Valid_Out & channel35_Kernel110_Valid_Out & channel36_Kernel110_Valid_Out & channel37_Kernel110_Valid_Out & channel38_Kernel110_Valid_Out & channel39_Kernel110_Valid_Out & channel40_Kernel110_Valid_Out & channel41_Kernel110_Valid_Out & channel42_Kernel110_Valid_Out & channel43_Kernel110_Valid_Out & channel44_Kernel110_Valid_Out & channel45_Kernel110_Valid_Out & channel46_Kernel110_Valid_Out & channel47_Kernel110_Valid_Out & channel48_Kernel110_Valid_Out & channel49_Kernel110_Valid_Out & channel50_Kernel110_Valid_Out & channel51_Kernel110_Valid_Out & channel52_Kernel110_Valid_Out & channel53_Kernel110_Valid_Out & channel54_Kernel110_Valid_Out & channel55_Kernel110_Valid_Out & channel56_Kernel110_Valid_Out & channel57_Kernel110_Valid_Out & channel58_Kernel110_Valid_Out & channel59_Kernel110_Valid_Out & channel60_Kernel110_Valid_Out & channel61_Kernel110_Valid_Out & channel62_Kernel110_Valid_Out & channel63_Kernel110_Valid_Out & channel64_Kernel110_Valid_Out;

	wire channel1_Kernel111_Valid_Out, channel2_Kernel111_Valid_Out, channel3_Kernel111_Valid_Out, channel4_Kernel111_Valid_Out, channel5_Kernel111_Valid_Out, channel6_Kernel111_Valid_Out, channel7_Kernel111_Valid_Out, channel8_Kernel111_Valid_Out, channel9_Kernel111_Valid_Out, channel10_Kernel111_Valid_Out, channel11_Kernel111_Valid_Out, channel12_Kernel111_Valid_Out, channel13_Kernel111_Valid_Out, channel14_Kernel111_Valid_Out, channel15_Kernel111_Valid_Out, channel16_Kernel111_Valid_Out, channel17_Kernel111_Valid_Out, channel18_Kernel111_Valid_Out, channel19_Kernel111_Valid_Out, channel20_Kernel111_Valid_Out, channel21_Kernel111_Valid_Out, channel22_Kernel111_Valid_Out, channel23_Kernel111_Valid_Out, channel24_Kernel111_Valid_Out, channel25_Kernel111_Valid_Out, channel26_Kernel111_Valid_Out, channel27_Kernel111_Valid_Out, channel28_Kernel111_Valid_Out, channel29_Kernel111_Valid_Out, channel30_Kernel111_Valid_Out, channel31_Kernel111_Valid_Out, channel32_Kernel111_Valid_Out, channel33_Kernel111_Valid_Out, channel34_Kernel111_Valid_Out, channel35_Kernel111_Valid_Out, channel36_Kernel111_Valid_Out, channel37_Kernel111_Valid_Out, channel38_Kernel111_Valid_Out, channel39_Kernel111_Valid_Out, channel40_Kernel111_Valid_Out, channel41_Kernel111_Valid_Out, channel42_Kernel111_Valid_Out, channel43_Kernel111_Valid_Out, channel44_Kernel111_Valid_Out, channel45_Kernel111_Valid_Out, channel46_Kernel111_Valid_Out, channel47_Kernel111_Valid_Out, channel48_Kernel111_Valid_Out, channel49_Kernel111_Valid_Out, channel50_Kernel111_Valid_Out, channel51_Kernel111_Valid_Out, channel52_Kernel111_Valid_Out, channel53_Kernel111_Valid_Out, channel54_Kernel111_Valid_Out, channel55_Kernel111_Valid_Out, channel56_Kernel111_Valid_Out, channel57_Kernel111_Valid_Out, channel58_Kernel111_Valid_Out, channel59_Kernel111_Valid_Out, channel60_Kernel111_Valid_Out, channel61_Kernel111_Valid_Out, channel62_Kernel111_Valid_Out, channel63_Kernel111_Valid_Out, channel64_Kernel111_Valid_Out;

	assign add_kernel111=channel1_Kernel111_Valid_Out & channel2_Kernel111_Valid_Out & channel3_Kernel111_Valid_Out & channel4_Kernel111_Valid_Out & channel5_Kernel111_Valid_Out & channel6_Kernel111_Valid_Out & channel7_Kernel111_Valid_Out & channel8_Kernel111_Valid_Out & channel9_Kernel111_Valid_Out & channel10_Kernel111_Valid_Out & channel11_Kernel111_Valid_Out & channel12_Kernel111_Valid_Out & channel13_Kernel111_Valid_Out & channel14_Kernel111_Valid_Out & channel15_Kernel111_Valid_Out & channel16_Kernel111_Valid_Out & channel17_Kernel111_Valid_Out & channel18_Kernel111_Valid_Out & channel19_Kernel111_Valid_Out & channel20_Kernel111_Valid_Out & channel21_Kernel111_Valid_Out & channel22_Kernel111_Valid_Out & channel23_Kernel111_Valid_Out & channel24_Kernel111_Valid_Out & channel25_Kernel111_Valid_Out & channel26_Kernel111_Valid_Out & channel27_Kernel111_Valid_Out & channel28_Kernel111_Valid_Out & channel29_Kernel111_Valid_Out & channel30_Kernel111_Valid_Out & channel31_Kernel111_Valid_Out & channel32_Kernel111_Valid_Out & channel33_Kernel111_Valid_Out & channel34_Kernel111_Valid_Out & channel35_Kernel111_Valid_Out & channel36_Kernel111_Valid_Out & channel37_Kernel111_Valid_Out & channel38_Kernel111_Valid_Out & channel39_Kernel111_Valid_Out & channel40_Kernel111_Valid_Out & channel41_Kernel111_Valid_Out & channel42_Kernel111_Valid_Out & channel43_Kernel111_Valid_Out & channel44_Kernel111_Valid_Out & channel45_Kernel111_Valid_Out & channel46_Kernel111_Valid_Out & channel47_Kernel111_Valid_Out & channel48_Kernel111_Valid_Out & channel49_Kernel111_Valid_Out & channel50_Kernel111_Valid_Out & channel51_Kernel111_Valid_Out & channel52_Kernel111_Valid_Out & channel53_Kernel111_Valid_Out & channel54_Kernel111_Valid_Out & channel55_Kernel111_Valid_Out & channel56_Kernel111_Valid_Out & channel57_Kernel111_Valid_Out & channel58_Kernel111_Valid_Out & channel59_Kernel111_Valid_Out & channel60_Kernel111_Valid_Out & channel61_Kernel111_Valid_Out & channel62_Kernel111_Valid_Out & channel63_Kernel111_Valid_Out & channel64_Kernel111_Valid_Out;

	wire channel1_Kernel112_Valid_Out, channel2_Kernel112_Valid_Out, channel3_Kernel112_Valid_Out, channel4_Kernel112_Valid_Out, channel5_Kernel112_Valid_Out, channel6_Kernel112_Valid_Out, channel7_Kernel112_Valid_Out, channel8_Kernel112_Valid_Out, channel9_Kernel112_Valid_Out, channel10_Kernel112_Valid_Out, channel11_Kernel112_Valid_Out, channel12_Kernel112_Valid_Out, channel13_Kernel112_Valid_Out, channel14_Kernel112_Valid_Out, channel15_Kernel112_Valid_Out, channel16_Kernel112_Valid_Out, channel17_Kernel112_Valid_Out, channel18_Kernel112_Valid_Out, channel19_Kernel112_Valid_Out, channel20_Kernel112_Valid_Out, channel21_Kernel112_Valid_Out, channel22_Kernel112_Valid_Out, channel23_Kernel112_Valid_Out, channel24_Kernel112_Valid_Out, channel25_Kernel112_Valid_Out, channel26_Kernel112_Valid_Out, channel27_Kernel112_Valid_Out, channel28_Kernel112_Valid_Out, channel29_Kernel112_Valid_Out, channel30_Kernel112_Valid_Out, channel31_Kernel112_Valid_Out, channel32_Kernel112_Valid_Out, channel33_Kernel112_Valid_Out, channel34_Kernel112_Valid_Out, channel35_Kernel112_Valid_Out, channel36_Kernel112_Valid_Out, channel37_Kernel112_Valid_Out, channel38_Kernel112_Valid_Out, channel39_Kernel112_Valid_Out, channel40_Kernel112_Valid_Out, channel41_Kernel112_Valid_Out, channel42_Kernel112_Valid_Out, channel43_Kernel112_Valid_Out, channel44_Kernel112_Valid_Out, channel45_Kernel112_Valid_Out, channel46_Kernel112_Valid_Out, channel47_Kernel112_Valid_Out, channel48_Kernel112_Valid_Out, channel49_Kernel112_Valid_Out, channel50_Kernel112_Valid_Out, channel51_Kernel112_Valid_Out, channel52_Kernel112_Valid_Out, channel53_Kernel112_Valid_Out, channel54_Kernel112_Valid_Out, channel55_Kernel112_Valid_Out, channel56_Kernel112_Valid_Out, channel57_Kernel112_Valid_Out, channel58_Kernel112_Valid_Out, channel59_Kernel112_Valid_Out, channel60_Kernel112_Valid_Out, channel61_Kernel112_Valid_Out, channel62_Kernel112_Valid_Out, channel63_Kernel112_Valid_Out, channel64_Kernel112_Valid_Out;

	assign add_kernel112=channel1_Kernel112_Valid_Out & channel2_Kernel112_Valid_Out & channel3_Kernel112_Valid_Out & channel4_Kernel112_Valid_Out & channel5_Kernel112_Valid_Out & channel6_Kernel112_Valid_Out & channel7_Kernel112_Valid_Out & channel8_Kernel112_Valid_Out & channel9_Kernel112_Valid_Out & channel10_Kernel112_Valid_Out & channel11_Kernel112_Valid_Out & channel12_Kernel112_Valid_Out & channel13_Kernel112_Valid_Out & channel14_Kernel112_Valid_Out & channel15_Kernel112_Valid_Out & channel16_Kernel112_Valid_Out & channel17_Kernel112_Valid_Out & channel18_Kernel112_Valid_Out & channel19_Kernel112_Valid_Out & channel20_Kernel112_Valid_Out & channel21_Kernel112_Valid_Out & channel22_Kernel112_Valid_Out & channel23_Kernel112_Valid_Out & channel24_Kernel112_Valid_Out & channel25_Kernel112_Valid_Out & channel26_Kernel112_Valid_Out & channel27_Kernel112_Valid_Out & channel28_Kernel112_Valid_Out & channel29_Kernel112_Valid_Out & channel30_Kernel112_Valid_Out & channel31_Kernel112_Valid_Out & channel32_Kernel112_Valid_Out & channel33_Kernel112_Valid_Out & channel34_Kernel112_Valid_Out & channel35_Kernel112_Valid_Out & channel36_Kernel112_Valid_Out & channel37_Kernel112_Valid_Out & channel38_Kernel112_Valid_Out & channel39_Kernel112_Valid_Out & channel40_Kernel112_Valid_Out & channel41_Kernel112_Valid_Out & channel42_Kernel112_Valid_Out & channel43_Kernel112_Valid_Out & channel44_Kernel112_Valid_Out & channel45_Kernel112_Valid_Out & channel46_Kernel112_Valid_Out & channel47_Kernel112_Valid_Out & channel48_Kernel112_Valid_Out & channel49_Kernel112_Valid_Out & channel50_Kernel112_Valid_Out & channel51_Kernel112_Valid_Out & channel52_Kernel112_Valid_Out & channel53_Kernel112_Valid_Out & channel54_Kernel112_Valid_Out & channel55_Kernel112_Valid_Out & channel56_Kernel112_Valid_Out & channel57_Kernel112_Valid_Out & channel58_Kernel112_Valid_Out & channel59_Kernel112_Valid_Out & channel60_Kernel112_Valid_Out & channel61_Kernel112_Valid_Out & channel62_Kernel112_Valid_Out & channel63_Kernel112_Valid_Out & channel64_Kernel112_Valid_Out;

	wire channel1_Kernel113_Valid_Out, channel2_Kernel113_Valid_Out, channel3_Kernel113_Valid_Out, channel4_Kernel113_Valid_Out, channel5_Kernel113_Valid_Out, channel6_Kernel113_Valid_Out, channel7_Kernel113_Valid_Out, channel8_Kernel113_Valid_Out, channel9_Kernel113_Valid_Out, channel10_Kernel113_Valid_Out, channel11_Kernel113_Valid_Out, channel12_Kernel113_Valid_Out, channel13_Kernel113_Valid_Out, channel14_Kernel113_Valid_Out, channel15_Kernel113_Valid_Out, channel16_Kernel113_Valid_Out, channel17_Kernel113_Valid_Out, channel18_Kernel113_Valid_Out, channel19_Kernel113_Valid_Out, channel20_Kernel113_Valid_Out, channel21_Kernel113_Valid_Out, channel22_Kernel113_Valid_Out, channel23_Kernel113_Valid_Out, channel24_Kernel113_Valid_Out, channel25_Kernel113_Valid_Out, channel26_Kernel113_Valid_Out, channel27_Kernel113_Valid_Out, channel28_Kernel113_Valid_Out, channel29_Kernel113_Valid_Out, channel30_Kernel113_Valid_Out, channel31_Kernel113_Valid_Out, channel32_Kernel113_Valid_Out, channel33_Kernel113_Valid_Out, channel34_Kernel113_Valid_Out, channel35_Kernel113_Valid_Out, channel36_Kernel113_Valid_Out, channel37_Kernel113_Valid_Out, channel38_Kernel113_Valid_Out, channel39_Kernel113_Valid_Out, channel40_Kernel113_Valid_Out, channel41_Kernel113_Valid_Out, channel42_Kernel113_Valid_Out, channel43_Kernel113_Valid_Out, channel44_Kernel113_Valid_Out, channel45_Kernel113_Valid_Out, channel46_Kernel113_Valid_Out, channel47_Kernel113_Valid_Out, channel48_Kernel113_Valid_Out, channel49_Kernel113_Valid_Out, channel50_Kernel113_Valid_Out, channel51_Kernel113_Valid_Out, channel52_Kernel113_Valid_Out, channel53_Kernel113_Valid_Out, channel54_Kernel113_Valid_Out, channel55_Kernel113_Valid_Out, channel56_Kernel113_Valid_Out, channel57_Kernel113_Valid_Out, channel58_Kernel113_Valid_Out, channel59_Kernel113_Valid_Out, channel60_Kernel113_Valid_Out, channel61_Kernel113_Valid_Out, channel62_Kernel113_Valid_Out, channel63_Kernel113_Valid_Out, channel64_Kernel113_Valid_Out;

	assign add_kernel113=channel1_Kernel113_Valid_Out & channel2_Kernel113_Valid_Out & channel3_Kernel113_Valid_Out & channel4_Kernel113_Valid_Out & channel5_Kernel113_Valid_Out & channel6_Kernel113_Valid_Out & channel7_Kernel113_Valid_Out & channel8_Kernel113_Valid_Out & channel9_Kernel113_Valid_Out & channel10_Kernel113_Valid_Out & channel11_Kernel113_Valid_Out & channel12_Kernel113_Valid_Out & channel13_Kernel113_Valid_Out & channel14_Kernel113_Valid_Out & channel15_Kernel113_Valid_Out & channel16_Kernel113_Valid_Out & channel17_Kernel113_Valid_Out & channel18_Kernel113_Valid_Out & channel19_Kernel113_Valid_Out & channel20_Kernel113_Valid_Out & channel21_Kernel113_Valid_Out & channel22_Kernel113_Valid_Out & channel23_Kernel113_Valid_Out & channel24_Kernel113_Valid_Out & channel25_Kernel113_Valid_Out & channel26_Kernel113_Valid_Out & channel27_Kernel113_Valid_Out & channel28_Kernel113_Valid_Out & channel29_Kernel113_Valid_Out & channel30_Kernel113_Valid_Out & channel31_Kernel113_Valid_Out & channel32_Kernel113_Valid_Out & channel33_Kernel113_Valid_Out & channel34_Kernel113_Valid_Out & channel35_Kernel113_Valid_Out & channel36_Kernel113_Valid_Out & channel37_Kernel113_Valid_Out & channel38_Kernel113_Valid_Out & channel39_Kernel113_Valid_Out & channel40_Kernel113_Valid_Out & channel41_Kernel113_Valid_Out & channel42_Kernel113_Valid_Out & channel43_Kernel113_Valid_Out & channel44_Kernel113_Valid_Out & channel45_Kernel113_Valid_Out & channel46_Kernel113_Valid_Out & channel47_Kernel113_Valid_Out & channel48_Kernel113_Valid_Out & channel49_Kernel113_Valid_Out & channel50_Kernel113_Valid_Out & channel51_Kernel113_Valid_Out & channel52_Kernel113_Valid_Out & channel53_Kernel113_Valid_Out & channel54_Kernel113_Valid_Out & channel55_Kernel113_Valid_Out & channel56_Kernel113_Valid_Out & channel57_Kernel113_Valid_Out & channel58_Kernel113_Valid_Out & channel59_Kernel113_Valid_Out & channel60_Kernel113_Valid_Out & channel61_Kernel113_Valid_Out & channel62_Kernel113_Valid_Out & channel63_Kernel113_Valid_Out & channel64_Kernel113_Valid_Out;

	wire channel1_Kernel114_Valid_Out, channel2_Kernel114_Valid_Out, channel3_Kernel114_Valid_Out, channel4_Kernel114_Valid_Out, channel5_Kernel114_Valid_Out, channel6_Kernel114_Valid_Out, channel7_Kernel114_Valid_Out, channel8_Kernel114_Valid_Out, channel9_Kernel114_Valid_Out, channel10_Kernel114_Valid_Out, channel11_Kernel114_Valid_Out, channel12_Kernel114_Valid_Out, channel13_Kernel114_Valid_Out, channel14_Kernel114_Valid_Out, channel15_Kernel114_Valid_Out, channel16_Kernel114_Valid_Out, channel17_Kernel114_Valid_Out, channel18_Kernel114_Valid_Out, channel19_Kernel114_Valid_Out, channel20_Kernel114_Valid_Out, channel21_Kernel114_Valid_Out, channel22_Kernel114_Valid_Out, channel23_Kernel114_Valid_Out, channel24_Kernel114_Valid_Out, channel25_Kernel114_Valid_Out, channel26_Kernel114_Valid_Out, channel27_Kernel114_Valid_Out, channel28_Kernel114_Valid_Out, channel29_Kernel114_Valid_Out, channel30_Kernel114_Valid_Out, channel31_Kernel114_Valid_Out, channel32_Kernel114_Valid_Out, channel33_Kernel114_Valid_Out, channel34_Kernel114_Valid_Out, channel35_Kernel114_Valid_Out, channel36_Kernel114_Valid_Out, channel37_Kernel114_Valid_Out, channel38_Kernel114_Valid_Out, channel39_Kernel114_Valid_Out, channel40_Kernel114_Valid_Out, channel41_Kernel114_Valid_Out, channel42_Kernel114_Valid_Out, channel43_Kernel114_Valid_Out, channel44_Kernel114_Valid_Out, channel45_Kernel114_Valid_Out, channel46_Kernel114_Valid_Out, channel47_Kernel114_Valid_Out, channel48_Kernel114_Valid_Out, channel49_Kernel114_Valid_Out, channel50_Kernel114_Valid_Out, channel51_Kernel114_Valid_Out, channel52_Kernel114_Valid_Out, channel53_Kernel114_Valid_Out, channel54_Kernel114_Valid_Out, channel55_Kernel114_Valid_Out, channel56_Kernel114_Valid_Out, channel57_Kernel114_Valid_Out, channel58_Kernel114_Valid_Out, channel59_Kernel114_Valid_Out, channel60_Kernel114_Valid_Out, channel61_Kernel114_Valid_Out, channel62_Kernel114_Valid_Out, channel63_Kernel114_Valid_Out, channel64_Kernel114_Valid_Out;

	assign add_kernel114=channel1_Kernel114_Valid_Out & channel2_Kernel114_Valid_Out & channel3_Kernel114_Valid_Out & channel4_Kernel114_Valid_Out & channel5_Kernel114_Valid_Out & channel6_Kernel114_Valid_Out & channel7_Kernel114_Valid_Out & channel8_Kernel114_Valid_Out & channel9_Kernel114_Valid_Out & channel10_Kernel114_Valid_Out & channel11_Kernel114_Valid_Out & channel12_Kernel114_Valid_Out & channel13_Kernel114_Valid_Out & channel14_Kernel114_Valid_Out & channel15_Kernel114_Valid_Out & channel16_Kernel114_Valid_Out & channel17_Kernel114_Valid_Out & channel18_Kernel114_Valid_Out & channel19_Kernel114_Valid_Out & channel20_Kernel114_Valid_Out & channel21_Kernel114_Valid_Out & channel22_Kernel114_Valid_Out & channel23_Kernel114_Valid_Out & channel24_Kernel114_Valid_Out & channel25_Kernel114_Valid_Out & channel26_Kernel114_Valid_Out & channel27_Kernel114_Valid_Out & channel28_Kernel114_Valid_Out & channel29_Kernel114_Valid_Out & channel30_Kernel114_Valid_Out & channel31_Kernel114_Valid_Out & channel32_Kernel114_Valid_Out & channel33_Kernel114_Valid_Out & channel34_Kernel114_Valid_Out & channel35_Kernel114_Valid_Out & channel36_Kernel114_Valid_Out & channel37_Kernel114_Valid_Out & channel38_Kernel114_Valid_Out & channel39_Kernel114_Valid_Out & channel40_Kernel114_Valid_Out & channel41_Kernel114_Valid_Out & channel42_Kernel114_Valid_Out & channel43_Kernel114_Valid_Out & channel44_Kernel114_Valid_Out & channel45_Kernel114_Valid_Out & channel46_Kernel114_Valid_Out & channel47_Kernel114_Valid_Out & channel48_Kernel114_Valid_Out & channel49_Kernel114_Valid_Out & channel50_Kernel114_Valid_Out & channel51_Kernel114_Valid_Out & channel52_Kernel114_Valid_Out & channel53_Kernel114_Valid_Out & channel54_Kernel114_Valid_Out & channel55_Kernel114_Valid_Out & channel56_Kernel114_Valid_Out & channel57_Kernel114_Valid_Out & channel58_Kernel114_Valid_Out & channel59_Kernel114_Valid_Out & channel60_Kernel114_Valid_Out & channel61_Kernel114_Valid_Out & channel62_Kernel114_Valid_Out & channel63_Kernel114_Valid_Out & channel64_Kernel114_Valid_Out;

	wire channel1_Kernel115_Valid_Out, channel2_Kernel115_Valid_Out, channel3_Kernel115_Valid_Out, channel4_Kernel115_Valid_Out, channel5_Kernel115_Valid_Out, channel6_Kernel115_Valid_Out, channel7_Kernel115_Valid_Out, channel8_Kernel115_Valid_Out, channel9_Kernel115_Valid_Out, channel10_Kernel115_Valid_Out, channel11_Kernel115_Valid_Out, channel12_Kernel115_Valid_Out, channel13_Kernel115_Valid_Out, channel14_Kernel115_Valid_Out, channel15_Kernel115_Valid_Out, channel16_Kernel115_Valid_Out, channel17_Kernel115_Valid_Out, channel18_Kernel115_Valid_Out, channel19_Kernel115_Valid_Out, channel20_Kernel115_Valid_Out, channel21_Kernel115_Valid_Out, channel22_Kernel115_Valid_Out, channel23_Kernel115_Valid_Out, channel24_Kernel115_Valid_Out, channel25_Kernel115_Valid_Out, channel26_Kernel115_Valid_Out, channel27_Kernel115_Valid_Out, channel28_Kernel115_Valid_Out, channel29_Kernel115_Valid_Out, channel30_Kernel115_Valid_Out, channel31_Kernel115_Valid_Out, channel32_Kernel115_Valid_Out, channel33_Kernel115_Valid_Out, channel34_Kernel115_Valid_Out, channel35_Kernel115_Valid_Out, channel36_Kernel115_Valid_Out, channel37_Kernel115_Valid_Out, channel38_Kernel115_Valid_Out, channel39_Kernel115_Valid_Out, channel40_Kernel115_Valid_Out, channel41_Kernel115_Valid_Out, channel42_Kernel115_Valid_Out, channel43_Kernel115_Valid_Out, channel44_Kernel115_Valid_Out, channel45_Kernel115_Valid_Out, channel46_Kernel115_Valid_Out, channel47_Kernel115_Valid_Out, channel48_Kernel115_Valid_Out, channel49_Kernel115_Valid_Out, channel50_Kernel115_Valid_Out, channel51_Kernel115_Valid_Out, channel52_Kernel115_Valid_Out, channel53_Kernel115_Valid_Out, channel54_Kernel115_Valid_Out, channel55_Kernel115_Valid_Out, channel56_Kernel115_Valid_Out, channel57_Kernel115_Valid_Out, channel58_Kernel115_Valid_Out, channel59_Kernel115_Valid_Out, channel60_Kernel115_Valid_Out, channel61_Kernel115_Valid_Out, channel62_Kernel115_Valid_Out, channel63_Kernel115_Valid_Out, channel64_Kernel115_Valid_Out;

	assign add_kernel115=channel1_Kernel115_Valid_Out & channel2_Kernel115_Valid_Out & channel3_Kernel115_Valid_Out & channel4_Kernel115_Valid_Out & channel5_Kernel115_Valid_Out & channel6_Kernel115_Valid_Out & channel7_Kernel115_Valid_Out & channel8_Kernel115_Valid_Out & channel9_Kernel115_Valid_Out & channel10_Kernel115_Valid_Out & channel11_Kernel115_Valid_Out & channel12_Kernel115_Valid_Out & channel13_Kernel115_Valid_Out & channel14_Kernel115_Valid_Out & channel15_Kernel115_Valid_Out & channel16_Kernel115_Valid_Out & channel17_Kernel115_Valid_Out & channel18_Kernel115_Valid_Out & channel19_Kernel115_Valid_Out & channel20_Kernel115_Valid_Out & channel21_Kernel115_Valid_Out & channel22_Kernel115_Valid_Out & channel23_Kernel115_Valid_Out & channel24_Kernel115_Valid_Out & channel25_Kernel115_Valid_Out & channel26_Kernel115_Valid_Out & channel27_Kernel115_Valid_Out & channel28_Kernel115_Valid_Out & channel29_Kernel115_Valid_Out & channel30_Kernel115_Valid_Out & channel31_Kernel115_Valid_Out & channel32_Kernel115_Valid_Out & channel33_Kernel115_Valid_Out & channel34_Kernel115_Valid_Out & channel35_Kernel115_Valid_Out & channel36_Kernel115_Valid_Out & channel37_Kernel115_Valid_Out & channel38_Kernel115_Valid_Out & channel39_Kernel115_Valid_Out & channel40_Kernel115_Valid_Out & channel41_Kernel115_Valid_Out & channel42_Kernel115_Valid_Out & channel43_Kernel115_Valid_Out & channel44_Kernel115_Valid_Out & channel45_Kernel115_Valid_Out & channel46_Kernel115_Valid_Out & channel47_Kernel115_Valid_Out & channel48_Kernel115_Valid_Out & channel49_Kernel115_Valid_Out & channel50_Kernel115_Valid_Out & channel51_Kernel115_Valid_Out & channel52_Kernel115_Valid_Out & channel53_Kernel115_Valid_Out & channel54_Kernel115_Valid_Out & channel55_Kernel115_Valid_Out & channel56_Kernel115_Valid_Out & channel57_Kernel115_Valid_Out & channel58_Kernel115_Valid_Out & channel59_Kernel115_Valid_Out & channel60_Kernel115_Valid_Out & channel61_Kernel115_Valid_Out & channel62_Kernel115_Valid_Out & channel63_Kernel115_Valid_Out & channel64_Kernel115_Valid_Out;

	wire channel1_Kernel116_Valid_Out, channel2_Kernel116_Valid_Out, channel3_Kernel116_Valid_Out, channel4_Kernel116_Valid_Out, channel5_Kernel116_Valid_Out, channel6_Kernel116_Valid_Out, channel7_Kernel116_Valid_Out, channel8_Kernel116_Valid_Out, channel9_Kernel116_Valid_Out, channel10_Kernel116_Valid_Out, channel11_Kernel116_Valid_Out, channel12_Kernel116_Valid_Out, channel13_Kernel116_Valid_Out, channel14_Kernel116_Valid_Out, channel15_Kernel116_Valid_Out, channel16_Kernel116_Valid_Out, channel17_Kernel116_Valid_Out, channel18_Kernel116_Valid_Out, channel19_Kernel116_Valid_Out, channel20_Kernel116_Valid_Out, channel21_Kernel116_Valid_Out, channel22_Kernel116_Valid_Out, channel23_Kernel116_Valid_Out, channel24_Kernel116_Valid_Out, channel25_Kernel116_Valid_Out, channel26_Kernel116_Valid_Out, channel27_Kernel116_Valid_Out, channel28_Kernel116_Valid_Out, channel29_Kernel116_Valid_Out, channel30_Kernel116_Valid_Out, channel31_Kernel116_Valid_Out, channel32_Kernel116_Valid_Out, channel33_Kernel116_Valid_Out, channel34_Kernel116_Valid_Out, channel35_Kernel116_Valid_Out, channel36_Kernel116_Valid_Out, channel37_Kernel116_Valid_Out, channel38_Kernel116_Valid_Out, channel39_Kernel116_Valid_Out, channel40_Kernel116_Valid_Out, channel41_Kernel116_Valid_Out, channel42_Kernel116_Valid_Out, channel43_Kernel116_Valid_Out, channel44_Kernel116_Valid_Out, channel45_Kernel116_Valid_Out, channel46_Kernel116_Valid_Out, channel47_Kernel116_Valid_Out, channel48_Kernel116_Valid_Out, channel49_Kernel116_Valid_Out, channel50_Kernel116_Valid_Out, channel51_Kernel116_Valid_Out, channel52_Kernel116_Valid_Out, channel53_Kernel116_Valid_Out, channel54_Kernel116_Valid_Out, channel55_Kernel116_Valid_Out, channel56_Kernel116_Valid_Out, channel57_Kernel116_Valid_Out, channel58_Kernel116_Valid_Out, channel59_Kernel116_Valid_Out, channel60_Kernel116_Valid_Out, channel61_Kernel116_Valid_Out, channel62_Kernel116_Valid_Out, channel63_Kernel116_Valid_Out, channel64_Kernel116_Valid_Out;

	assign add_kernel116=channel1_Kernel116_Valid_Out & channel2_Kernel116_Valid_Out & channel3_Kernel116_Valid_Out & channel4_Kernel116_Valid_Out & channel5_Kernel116_Valid_Out & channel6_Kernel116_Valid_Out & channel7_Kernel116_Valid_Out & channel8_Kernel116_Valid_Out & channel9_Kernel116_Valid_Out & channel10_Kernel116_Valid_Out & channel11_Kernel116_Valid_Out & channel12_Kernel116_Valid_Out & channel13_Kernel116_Valid_Out & channel14_Kernel116_Valid_Out & channel15_Kernel116_Valid_Out & channel16_Kernel116_Valid_Out & channel17_Kernel116_Valid_Out & channel18_Kernel116_Valid_Out & channel19_Kernel116_Valid_Out & channel20_Kernel116_Valid_Out & channel21_Kernel116_Valid_Out & channel22_Kernel116_Valid_Out & channel23_Kernel116_Valid_Out & channel24_Kernel116_Valid_Out & channel25_Kernel116_Valid_Out & channel26_Kernel116_Valid_Out & channel27_Kernel116_Valid_Out & channel28_Kernel116_Valid_Out & channel29_Kernel116_Valid_Out & channel30_Kernel116_Valid_Out & channel31_Kernel116_Valid_Out & channel32_Kernel116_Valid_Out & channel33_Kernel116_Valid_Out & channel34_Kernel116_Valid_Out & channel35_Kernel116_Valid_Out & channel36_Kernel116_Valid_Out & channel37_Kernel116_Valid_Out & channel38_Kernel116_Valid_Out & channel39_Kernel116_Valid_Out & channel40_Kernel116_Valid_Out & channel41_Kernel116_Valid_Out & channel42_Kernel116_Valid_Out & channel43_Kernel116_Valid_Out & channel44_Kernel116_Valid_Out & channel45_Kernel116_Valid_Out & channel46_Kernel116_Valid_Out & channel47_Kernel116_Valid_Out & channel48_Kernel116_Valid_Out & channel49_Kernel116_Valid_Out & channel50_Kernel116_Valid_Out & channel51_Kernel116_Valid_Out & channel52_Kernel116_Valid_Out & channel53_Kernel116_Valid_Out & channel54_Kernel116_Valid_Out & channel55_Kernel116_Valid_Out & channel56_Kernel116_Valid_Out & channel57_Kernel116_Valid_Out & channel58_Kernel116_Valid_Out & channel59_Kernel116_Valid_Out & channel60_Kernel116_Valid_Out & channel61_Kernel116_Valid_Out & channel62_Kernel116_Valid_Out & channel63_Kernel116_Valid_Out & channel64_Kernel116_Valid_Out;

	wire channel1_Kernel117_Valid_Out, channel2_Kernel117_Valid_Out, channel3_Kernel117_Valid_Out, channel4_Kernel117_Valid_Out, channel5_Kernel117_Valid_Out, channel6_Kernel117_Valid_Out, channel7_Kernel117_Valid_Out, channel8_Kernel117_Valid_Out, channel9_Kernel117_Valid_Out, channel10_Kernel117_Valid_Out, channel11_Kernel117_Valid_Out, channel12_Kernel117_Valid_Out, channel13_Kernel117_Valid_Out, channel14_Kernel117_Valid_Out, channel15_Kernel117_Valid_Out, channel16_Kernel117_Valid_Out, channel17_Kernel117_Valid_Out, channel18_Kernel117_Valid_Out, channel19_Kernel117_Valid_Out, channel20_Kernel117_Valid_Out, channel21_Kernel117_Valid_Out, channel22_Kernel117_Valid_Out, channel23_Kernel117_Valid_Out, channel24_Kernel117_Valid_Out, channel25_Kernel117_Valid_Out, channel26_Kernel117_Valid_Out, channel27_Kernel117_Valid_Out, channel28_Kernel117_Valid_Out, channel29_Kernel117_Valid_Out, channel30_Kernel117_Valid_Out, channel31_Kernel117_Valid_Out, channel32_Kernel117_Valid_Out, channel33_Kernel117_Valid_Out, channel34_Kernel117_Valid_Out, channel35_Kernel117_Valid_Out, channel36_Kernel117_Valid_Out, channel37_Kernel117_Valid_Out, channel38_Kernel117_Valid_Out, channel39_Kernel117_Valid_Out, channel40_Kernel117_Valid_Out, channel41_Kernel117_Valid_Out, channel42_Kernel117_Valid_Out, channel43_Kernel117_Valid_Out, channel44_Kernel117_Valid_Out, channel45_Kernel117_Valid_Out, channel46_Kernel117_Valid_Out, channel47_Kernel117_Valid_Out, channel48_Kernel117_Valid_Out, channel49_Kernel117_Valid_Out, channel50_Kernel117_Valid_Out, channel51_Kernel117_Valid_Out, channel52_Kernel117_Valid_Out, channel53_Kernel117_Valid_Out, channel54_Kernel117_Valid_Out, channel55_Kernel117_Valid_Out, channel56_Kernel117_Valid_Out, channel57_Kernel117_Valid_Out, channel58_Kernel117_Valid_Out, channel59_Kernel117_Valid_Out, channel60_Kernel117_Valid_Out, channel61_Kernel117_Valid_Out, channel62_Kernel117_Valid_Out, channel63_Kernel117_Valid_Out, channel64_Kernel117_Valid_Out;

	assign add_kernel117=channel1_Kernel117_Valid_Out & channel2_Kernel117_Valid_Out & channel3_Kernel117_Valid_Out & channel4_Kernel117_Valid_Out & channel5_Kernel117_Valid_Out & channel6_Kernel117_Valid_Out & channel7_Kernel117_Valid_Out & channel8_Kernel117_Valid_Out & channel9_Kernel117_Valid_Out & channel10_Kernel117_Valid_Out & channel11_Kernel117_Valid_Out & channel12_Kernel117_Valid_Out & channel13_Kernel117_Valid_Out & channel14_Kernel117_Valid_Out & channel15_Kernel117_Valid_Out & channel16_Kernel117_Valid_Out & channel17_Kernel117_Valid_Out & channel18_Kernel117_Valid_Out & channel19_Kernel117_Valid_Out & channel20_Kernel117_Valid_Out & channel21_Kernel117_Valid_Out & channel22_Kernel117_Valid_Out & channel23_Kernel117_Valid_Out & channel24_Kernel117_Valid_Out & channel25_Kernel117_Valid_Out & channel26_Kernel117_Valid_Out & channel27_Kernel117_Valid_Out & channel28_Kernel117_Valid_Out & channel29_Kernel117_Valid_Out & channel30_Kernel117_Valid_Out & channel31_Kernel117_Valid_Out & channel32_Kernel117_Valid_Out & channel33_Kernel117_Valid_Out & channel34_Kernel117_Valid_Out & channel35_Kernel117_Valid_Out & channel36_Kernel117_Valid_Out & channel37_Kernel117_Valid_Out & channel38_Kernel117_Valid_Out & channel39_Kernel117_Valid_Out & channel40_Kernel117_Valid_Out & channel41_Kernel117_Valid_Out & channel42_Kernel117_Valid_Out & channel43_Kernel117_Valid_Out & channel44_Kernel117_Valid_Out & channel45_Kernel117_Valid_Out & channel46_Kernel117_Valid_Out & channel47_Kernel117_Valid_Out & channel48_Kernel117_Valid_Out & channel49_Kernel117_Valid_Out & channel50_Kernel117_Valid_Out & channel51_Kernel117_Valid_Out & channel52_Kernel117_Valid_Out & channel53_Kernel117_Valid_Out & channel54_Kernel117_Valid_Out & channel55_Kernel117_Valid_Out & channel56_Kernel117_Valid_Out & channel57_Kernel117_Valid_Out & channel58_Kernel117_Valid_Out & channel59_Kernel117_Valid_Out & channel60_Kernel117_Valid_Out & channel61_Kernel117_Valid_Out & channel62_Kernel117_Valid_Out & channel63_Kernel117_Valid_Out & channel64_Kernel117_Valid_Out;

	wire channel1_Kernel118_Valid_Out, channel2_Kernel118_Valid_Out, channel3_Kernel118_Valid_Out, channel4_Kernel118_Valid_Out, channel5_Kernel118_Valid_Out, channel6_Kernel118_Valid_Out, channel7_Kernel118_Valid_Out, channel8_Kernel118_Valid_Out, channel9_Kernel118_Valid_Out, channel10_Kernel118_Valid_Out, channel11_Kernel118_Valid_Out, channel12_Kernel118_Valid_Out, channel13_Kernel118_Valid_Out, channel14_Kernel118_Valid_Out, channel15_Kernel118_Valid_Out, channel16_Kernel118_Valid_Out, channel17_Kernel118_Valid_Out, channel18_Kernel118_Valid_Out, channel19_Kernel118_Valid_Out, channel20_Kernel118_Valid_Out, channel21_Kernel118_Valid_Out, channel22_Kernel118_Valid_Out, channel23_Kernel118_Valid_Out, channel24_Kernel118_Valid_Out, channel25_Kernel118_Valid_Out, channel26_Kernel118_Valid_Out, channel27_Kernel118_Valid_Out, channel28_Kernel118_Valid_Out, channel29_Kernel118_Valid_Out, channel30_Kernel118_Valid_Out, channel31_Kernel118_Valid_Out, channel32_Kernel118_Valid_Out, channel33_Kernel118_Valid_Out, channel34_Kernel118_Valid_Out, channel35_Kernel118_Valid_Out, channel36_Kernel118_Valid_Out, channel37_Kernel118_Valid_Out, channel38_Kernel118_Valid_Out, channel39_Kernel118_Valid_Out, channel40_Kernel118_Valid_Out, channel41_Kernel118_Valid_Out, channel42_Kernel118_Valid_Out, channel43_Kernel118_Valid_Out, channel44_Kernel118_Valid_Out, channel45_Kernel118_Valid_Out, channel46_Kernel118_Valid_Out, channel47_Kernel118_Valid_Out, channel48_Kernel118_Valid_Out, channel49_Kernel118_Valid_Out, channel50_Kernel118_Valid_Out, channel51_Kernel118_Valid_Out, channel52_Kernel118_Valid_Out, channel53_Kernel118_Valid_Out, channel54_Kernel118_Valid_Out, channel55_Kernel118_Valid_Out, channel56_Kernel118_Valid_Out, channel57_Kernel118_Valid_Out, channel58_Kernel118_Valid_Out, channel59_Kernel118_Valid_Out, channel60_Kernel118_Valid_Out, channel61_Kernel118_Valid_Out, channel62_Kernel118_Valid_Out, channel63_Kernel118_Valid_Out, channel64_Kernel118_Valid_Out;

	assign add_kernel118=channel1_Kernel118_Valid_Out & channel2_Kernel118_Valid_Out & channel3_Kernel118_Valid_Out & channel4_Kernel118_Valid_Out & channel5_Kernel118_Valid_Out & channel6_Kernel118_Valid_Out & channel7_Kernel118_Valid_Out & channel8_Kernel118_Valid_Out & channel9_Kernel118_Valid_Out & channel10_Kernel118_Valid_Out & channel11_Kernel118_Valid_Out & channel12_Kernel118_Valid_Out & channel13_Kernel118_Valid_Out & channel14_Kernel118_Valid_Out & channel15_Kernel118_Valid_Out & channel16_Kernel118_Valid_Out & channel17_Kernel118_Valid_Out & channel18_Kernel118_Valid_Out & channel19_Kernel118_Valid_Out & channel20_Kernel118_Valid_Out & channel21_Kernel118_Valid_Out & channel22_Kernel118_Valid_Out & channel23_Kernel118_Valid_Out & channel24_Kernel118_Valid_Out & channel25_Kernel118_Valid_Out & channel26_Kernel118_Valid_Out & channel27_Kernel118_Valid_Out & channel28_Kernel118_Valid_Out & channel29_Kernel118_Valid_Out & channel30_Kernel118_Valid_Out & channel31_Kernel118_Valid_Out & channel32_Kernel118_Valid_Out & channel33_Kernel118_Valid_Out & channel34_Kernel118_Valid_Out & channel35_Kernel118_Valid_Out & channel36_Kernel118_Valid_Out & channel37_Kernel118_Valid_Out & channel38_Kernel118_Valid_Out & channel39_Kernel118_Valid_Out & channel40_Kernel118_Valid_Out & channel41_Kernel118_Valid_Out & channel42_Kernel118_Valid_Out & channel43_Kernel118_Valid_Out & channel44_Kernel118_Valid_Out & channel45_Kernel118_Valid_Out & channel46_Kernel118_Valid_Out & channel47_Kernel118_Valid_Out & channel48_Kernel118_Valid_Out & channel49_Kernel118_Valid_Out & channel50_Kernel118_Valid_Out & channel51_Kernel118_Valid_Out & channel52_Kernel118_Valid_Out & channel53_Kernel118_Valid_Out & channel54_Kernel118_Valid_Out & channel55_Kernel118_Valid_Out & channel56_Kernel118_Valid_Out & channel57_Kernel118_Valid_Out & channel58_Kernel118_Valid_Out & channel59_Kernel118_Valid_Out & channel60_Kernel118_Valid_Out & channel61_Kernel118_Valid_Out & channel62_Kernel118_Valid_Out & channel63_Kernel118_Valid_Out & channel64_Kernel118_Valid_Out;

	wire channel1_Kernel119_Valid_Out, channel2_Kernel119_Valid_Out, channel3_Kernel119_Valid_Out, channel4_Kernel119_Valid_Out, channel5_Kernel119_Valid_Out, channel6_Kernel119_Valid_Out, channel7_Kernel119_Valid_Out, channel8_Kernel119_Valid_Out, channel9_Kernel119_Valid_Out, channel10_Kernel119_Valid_Out, channel11_Kernel119_Valid_Out, channel12_Kernel119_Valid_Out, channel13_Kernel119_Valid_Out, channel14_Kernel119_Valid_Out, channel15_Kernel119_Valid_Out, channel16_Kernel119_Valid_Out, channel17_Kernel119_Valid_Out, channel18_Kernel119_Valid_Out, channel19_Kernel119_Valid_Out, channel20_Kernel119_Valid_Out, channel21_Kernel119_Valid_Out, channel22_Kernel119_Valid_Out, channel23_Kernel119_Valid_Out, channel24_Kernel119_Valid_Out, channel25_Kernel119_Valid_Out, channel26_Kernel119_Valid_Out, channel27_Kernel119_Valid_Out, channel28_Kernel119_Valid_Out, channel29_Kernel119_Valid_Out, channel30_Kernel119_Valid_Out, channel31_Kernel119_Valid_Out, channel32_Kernel119_Valid_Out, channel33_Kernel119_Valid_Out, channel34_Kernel119_Valid_Out, channel35_Kernel119_Valid_Out, channel36_Kernel119_Valid_Out, channel37_Kernel119_Valid_Out, channel38_Kernel119_Valid_Out, channel39_Kernel119_Valid_Out, channel40_Kernel119_Valid_Out, channel41_Kernel119_Valid_Out, channel42_Kernel119_Valid_Out, channel43_Kernel119_Valid_Out, channel44_Kernel119_Valid_Out, channel45_Kernel119_Valid_Out, channel46_Kernel119_Valid_Out, channel47_Kernel119_Valid_Out, channel48_Kernel119_Valid_Out, channel49_Kernel119_Valid_Out, channel50_Kernel119_Valid_Out, channel51_Kernel119_Valid_Out, channel52_Kernel119_Valid_Out, channel53_Kernel119_Valid_Out, channel54_Kernel119_Valid_Out, channel55_Kernel119_Valid_Out, channel56_Kernel119_Valid_Out, channel57_Kernel119_Valid_Out, channel58_Kernel119_Valid_Out, channel59_Kernel119_Valid_Out, channel60_Kernel119_Valid_Out, channel61_Kernel119_Valid_Out, channel62_Kernel119_Valid_Out, channel63_Kernel119_Valid_Out, channel64_Kernel119_Valid_Out;

	assign add_kernel119=channel1_Kernel119_Valid_Out & channel2_Kernel119_Valid_Out & channel3_Kernel119_Valid_Out & channel4_Kernel119_Valid_Out & channel5_Kernel119_Valid_Out & channel6_Kernel119_Valid_Out & channel7_Kernel119_Valid_Out & channel8_Kernel119_Valid_Out & channel9_Kernel119_Valid_Out & channel10_Kernel119_Valid_Out & channel11_Kernel119_Valid_Out & channel12_Kernel119_Valid_Out & channel13_Kernel119_Valid_Out & channel14_Kernel119_Valid_Out & channel15_Kernel119_Valid_Out & channel16_Kernel119_Valid_Out & channel17_Kernel119_Valid_Out & channel18_Kernel119_Valid_Out & channel19_Kernel119_Valid_Out & channel20_Kernel119_Valid_Out & channel21_Kernel119_Valid_Out & channel22_Kernel119_Valid_Out & channel23_Kernel119_Valid_Out & channel24_Kernel119_Valid_Out & channel25_Kernel119_Valid_Out & channel26_Kernel119_Valid_Out & channel27_Kernel119_Valid_Out & channel28_Kernel119_Valid_Out & channel29_Kernel119_Valid_Out & channel30_Kernel119_Valid_Out & channel31_Kernel119_Valid_Out & channel32_Kernel119_Valid_Out & channel33_Kernel119_Valid_Out & channel34_Kernel119_Valid_Out & channel35_Kernel119_Valid_Out & channel36_Kernel119_Valid_Out & channel37_Kernel119_Valid_Out & channel38_Kernel119_Valid_Out & channel39_Kernel119_Valid_Out & channel40_Kernel119_Valid_Out & channel41_Kernel119_Valid_Out & channel42_Kernel119_Valid_Out & channel43_Kernel119_Valid_Out & channel44_Kernel119_Valid_Out & channel45_Kernel119_Valid_Out & channel46_Kernel119_Valid_Out & channel47_Kernel119_Valid_Out & channel48_Kernel119_Valid_Out & channel49_Kernel119_Valid_Out & channel50_Kernel119_Valid_Out & channel51_Kernel119_Valid_Out & channel52_Kernel119_Valid_Out & channel53_Kernel119_Valid_Out & channel54_Kernel119_Valid_Out & channel55_Kernel119_Valid_Out & channel56_Kernel119_Valid_Out & channel57_Kernel119_Valid_Out & channel58_Kernel119_Valid_Out & channel59_Kernel119_Valid_Out & channel60_Kernel119_Valid_Out & channel61_Kernel119_Valid_Out & channel62_Kernel119_Valid_Out & channel63_Kernel119_Valid_Out & channel64_Kernel119_Valid_Out;

	wire channel1_Kernel120_Valid_Out, channel2_Kernel120_Valid_Out, channel3_Kernel120_Valid_Out, channel4_Kernel120_Valid_Out, channel5_Kernel120_Valid_Out, channel6_Kernel120_Valid_Out, channel7_Kernel120_Valid_Out, channel8_Kernel120_Valid_Out, channel9_Kernel120_Valid_Out, channel10_Kernel120_Valid_Out, channel11_Kernel120_Valid_Out, channel12_Kernel120_Valid_Out, channel13_Kernel120_Valid_Out, channel14_Kernel120_Valid_Out, channel15_Kernel120_Valid_Out, channel16_Kernel120_Valid_Out, channel17_Kernel120_Valid_Out, channel18_Kernel120_Valid_Out, channel19_Kernel120_Valid_Out, channel20_Kernel120_Valid_Out, channel21_Kernel120_Valid_Out, channel22_Kernel120_Valid_Out, channel23_Kernel120_Valid_Out, channel24_Kernel120_Valid_Out, channel25_Kernel120_Valid_Out, channel26_Kernel120_Valid_Out, channel27_Kernel120_Valid_Out, channel28_Kernel120_Valid_Out, channel29_Kernel120_Valid_Out, channel30_Kernel120_Valid_Out, channel31_Kernel120_Valid_Out, channel32_Kernel120_Valid_Out, channel33_Kernel120_Valid_Out, channel34_Kernel120_Valid_Out, channel35_Kernel120_Valid_Out, channel36_Kernel120_Valid_Out, channel37_Kernel120_Valid_Out, channel38_Kernel120_Valid_Out, channel39_Kernel120_Valid_Out, channel40_Kernel120_Valid_Out, channel41_Kernel120_Valid_Out, channel42_Kernel120_Valid_Out, channel43_Kernel120_Valid_Out, channel44_Kernel120_Valid_Out, channel45_Kernel120_Valid_Out, channel46_Kernel120_Valid_Out, channel47_Kernel120_Valid_Out, channel48_Kernel120_Valid_Out, channel49_Kernel120_Valid_Out, channel50_Kernel120_Valid_Out, channel51_Kernel120_Valid_Out, channel52_Kernel120_Valid_Out, channel53_Kernel120_Valid_Out, channel54_Kernel120_Valid_Out, channel55_Kernel120_Valid_Out, channel56_Kernel120_Valid_Out, channel57_Kernel120_Valid_Out, channel58_Kernel120_Valid_Out, channel59_Kernel120_Valid_Out, channel60_Kernel120_Valid_Out, channel61_Kernel120_Valid_Out, channel62_Kernel120_Valid_Out, channel63_Kernel120_Valid_Out, channel64_Kernel120_Valid_Out;

	assign add_kernel120=channel1_Kernel120_Valid_Out & channel2_Kernel120_Valid_Out & channel3_Kernel120_Valid_Out & channel4_Kernel120_Valid_Out & channel5_Kernel120_Valid_Out & channel6_Kernel120_Valid_Out & channel7_Kernel120_Valid_Out & channel8_Kernel120_Valid_Out & channel9_Kernel120_Valid_Out & channel10_Kernel120_Valid_Out & channel11_Kernel120_Valid_Out & channel12_Kernel120_Valid_Out & channel13_Kernel120_Valid_Out & channel14_Kernel120_Valid_Out & channel15_Kernel120_Valid_Out & channel16_Kernel120_Valid_Out & channel17_Kernel120_Valid_Out & channel18_Kernel120_Valid_Out & channel19_Kernel120_Valid_Out & channel20_Kernel120_Valid_Out & channel21_Kernel120_Valid_Out & channel22_Kernel120_Valid_Out & channel23_Kernel120_Valid_Out & channel24_Kernel120_Valid_Out & channel25_Kernel120_Valid_Out & channel26_Kernel120_Valid_Out & channel27_Kernel120_Valid_Out & channel28_Kernel120_Valid_Out & channel29_Kernel120_Valid_Out & channel30_Kernel120_Valid_Out & channel31_Kernel120_Valid_Out & channel32_Kernel120_Valid_Out & channel33_Kernel120_Valid_Out & channel34_Kernel120_Valid_Out & channel35_Kernel120_Valid_Out & channel36_Kernel120_Valid_Out & channel37_Kernel120_Valid_Out & channel38_Kernel120_Valid_Out & channel39_Kernel120_Valid_Out & channel40_Kernel120_Valid_Out & channel41_Kernel120_Valid_Out & channel42_Kernel120_Valid_Out & channel43_Kernel120_Valid_Out & channel44_Kernel120_Valid_Out & channel45_Kernel120_Valid_Out & channel46_Kernel120_Valid_Out & channel47_Kernel120_Valid_Out & channel48_Kernel120_Valid_Out & channel49_Kernel120_Valid_Out & channel50_Kernel120_Valid_Out & channel51_Kernel120_Valid_Out & channel52_Kernel120_Valid_Out & channel53_Kernel120_Valid_Out & channel54_Kernel120_Valid_Out & channel55_Kernel120_Valid_Out & channel56_Kernel120_Valid_Out & channel57_Kernel120_Valid_Out & channel58_Kernel120_Valid_Out & channel59_Kernel120_Valid_Out & channel60_Kernel120_Valid_Out & channel61_Kernel120_Valid_Out & channel62_Kernel120_Valid_Out & channel63_Kernel120_Valid_Out & channel64_Kernel120_Valid_Out;

	wire channel1_Kernel121_Valid_Out, channel2_Kernel121_Valid_Out, channel3_Kernel121_Valid_Out, channel4_Kernel121_Valid_Out, channel5_Kernel121_Valid_Out, channel6_Kernel121_Valid_Out, channel7_Kernel121_Valid_Out, channel8_Kernel121_Valid_Out, channel9_Kernel121_Valid_Out, channel10_Kernel121_Valid_Out, channel11_Kernel121_Valid_Out, channel12_Kernel121_Valid_Out, channel13_Kernel121_Valid_Out, channel14_Kernel121_Valid_Out, channel15_Kernel121_Valid_Out, channel16_Kernel121_Valid_Out, channel17_Kernel121_Valid_Out, channel18_Kernel121_Valid_Out, channel19_Kernel121_Valid_Out, channel20_Kernel121_Valid_Out, channel21_Kernel121_Valid_Out, channel22_Kernel121_Valid_Out, channel23_Kernel121_Valid_Out, channel24_Kernel121_Valid_Out, channel25_Kernel121_Valid_Out, channel26_Kernel121_Valid_Out, channel27_Kernel121_Valid_Out, channel28_Kernel121_Valid_Out, channel29_Kernel121_Valid_Out, channel30_Kernel121_Valid_Out, channel31_Kernel121_Valid_Out, channel32_Kernel121_Valid_Out, channel33_Kernel121_Valid_Out, channel34_Kernel121_Valid_Out, channel35_Kernel121_Valid_Out, channel36_Kernel121_Valid_Out, channel37_Kernel121_Valid_Out, channel38_Kernel121_Valid_Out, channel39_Kernel121_Valid_Out, channel40_Kernel121_Valid_Out, channel41_Kernel121_Valid_Out, channel42_Kernel121_Valid_Out, channel43_Kernel121_Valid_Out, channel44_Kernel121_Valid_Out, channel45_Kernel121_Valid_Out, channel46_Kernel121_Valid_Out, channel47_Kernel121_Valid_Out, channel48_Kernel121_Valid_Out, channel49_Kernel121_Valid_Out, channel50_Kernel121_Valid_Out, channel51_Kernel121_Valid_Out, channel52_Kernel121_Valid_Out, channel53_Kernel121_Valid_Out, channel54_Kernel121_Valid_Out, channel55_Kernel121_Valid_Out, channel56_Kernel121_Valid_Out, channel57_Kernel121_Valid_Out, channel58_Kernel121_Valid_Out, channel59_Kernel121_Valid_Out, channel60_Kernel121_Valid_Out, channel61_Kernel121_Valid_Out, channel62_Kernel121_Valid_Out, channel63_Kernel121_Valid_Out, channel64_Kernel121_Valid_Out;

	assign add_kernel121=channel1_Kernel121_Valid_Out & channel2_Kernel121_Valid_Out & channel3_Kernel121_Valid_Out & channel4_Kernel121_Valid_Out & channel5_Kernel121_Valid_Out & channel6_Kernel121_Valid_Out & channel7_Kernel121_Valid_Out & channel8_Kernel121_Valid_Out & channel9_Kernel121_Valid_Out & channel10_Kernel121_Valid_Out & channel11_Kernel121_Valid_Out & channel12_Kernel121_Valid_Out & channel13_Kernel121_Valid_Out & channel14_Kernel121_Valid_Out & channel15_Kernel121_Valid_Out & channel16_Kernel121_Valid_Out & channel17_Kernel121_Valid_Out & channel18_Kernel121_Valid_Out & channel19_Kernel121_Valid_Out & channel20_Kernel121_Valid_Out & channel21_Kernel121_Valid_Out & channel22_Kernel121_Valid_Out & channel23_Kernel121_Valid_Out & channel24_Kernel121_Valid_Out & channel25_Kernel121_Valid_Out & channel26_Kernel121_Valid_Out & channel27_Kernel121_Valid_Out & channel28_Kernel121_Valid_Out & channel29_Kernel121_Valid_Out & channel30_Kernel121_Valid_Out & channel31_Kernel121_Valid_Out & channel32_Kernel121_Valid_Out & channel33_Kernel121_Valid_Out & channel34_Kernel121_Valid_Out & channel35_Kernel121_Valid_Out & channel36_Kernel121_Valid_Out & channel37_Kernel121_Valid_Out & channel38_Kernel121_Valid_Out & channel39_Kernel121_Valid_Out & channel40_Kernel121_Valid_Out & channel41_Kernel121_Valid_Out & channel42_Kernel121_Valid_Out & channel43_Kernel121_Valid_Out & channel44_Kernel121_Valid_Out & channel45_Kernel121_Valid_Out & channel46_Kernel121_Valid_Out & channel47_Kernel121_Valid_Out & channel48_Kernel121_Valid_Out & channel49_Kernel121_Valid_Out & channel50_Kernel121_Valid_Out & channel51_Kernel121_Valid_Out & channel52_Kernel121_Valid_Out & channel53_Kernel121_Valid_Out & channel54_Kernel121_Valid_Out & channel55_Kernel121_Valid_Out & channel56_Kernel121_Valid_Out & channel57_Kernel121_Valid_Out & channel58_Kernel121_Valid_Out & channel59_Kernel121_Valid_Out & channel60_Kernel121_Valid_Out & channel61_Kernel121_Valid_Out & channel62_Kernel121_Valid_Out & channel63_Kernel121_Valid_Out & channel64_Kernel121_Valid_Out;

	wire channel1_Kernel122_Valid_Out, channel2_Kernel122_Valid_Out, channel3_Kernel122_Valid_Out, channel4_Kernel122_Valid_Out, channel5_Kernel122_Valid_Out, channel6_Kernel122_Valid_Out, channel7_Kernel122_Valid_Out, channel8_Kernel122_Valid_Out, channel9_Kernel122_Valid_Out, channel10_Kernel122_Valid_Out, channel11_Kernel122_Valid_Out, channel12_Kernel122_Valid_Out, channel13_Kernel122_Valid_Out, channel14_Kernel122_Valid_Out, channel15_Kernel122_Valid_Out, channel16_Kernel122_Valid_Out, channel17_Kernel122_Valid_Out, channel18_Kernel122_Valid_Out, channel19_Kernel122_Valid_Out, channel20_Kernel122_Valid_Out, channel21_Kernel122_Valid_Out, channel22_Kernel122_Valid_Out, channel23_Kernel122_Valid_Out, channel24_Kernel122_Valid_Out, channel25_Kernel122_Valid_Out, channel26_Kernel122_Valid_Out, channel27_Kernel122_Valid_Out, channel28_Kernel122_Valid_Out, channel29_Kernel122_Valid_Out, channel30_Kernel122_Valid_Out, channel31_Kernel122_Valid_Out, channel32_Kernel122_Valid_Out, channel33_Kernel122_Valid_Out, channel34_Kernel122_Valid_Out, channel35_Kernel122_Valid_Out, channel36_Kernel122_Valid_Out, channel37_Kernel122_Valid_Out, channel38_Kernel122_Valid_Out, channel39_Kernel122_Valid_Out, channel40_Kernel122_Valid_Out, channel41_Kernel122_Valid_Out, channel42_Kernel122_Valid_Out, channel43_Kernel122_Valid_Out, channel44_Kernel122_Valid_Out, channel45_Kernel122_Valid_Out, channel46_Kernel122_Valid_Out, channel47_Kernel122_Valid_Out, channel48_Kernel122_Valid_Out, channel49_Kernel122_Valid_Out, channel50_Kernel122_Valid_Out, channel51_Kernel122_Valid_Out, channel52_Kernel122_Valid_Out, channel53_Kernel122_Valid_Out, channel54_Kernel122_Valid_Out, channel55_Kernel122_Valid_Out, channel56_Kernel122_Valid_Out, channel57_Kernel122_Valid_Out, channel58_Kernel122_Valid_Out, channel59_Kernel122_Valid_Out, channel60_Kernel122_Valid_Out, channel61_Kernel122_Valid_Out, channel62_Kernel122_Valid_Out, channel63_Kernel122_Valid_Out, channel64_Kernel122_Valid_Out;

	assign add_kernel122=channel1_Kernel122_Valid_Out & channel2_Kernel122_Valid_Out & channel3_Kernel122_Valid_Out & channel4_Kernel122_Valid_Out & channel5_Kernel122_Valid_Out & channel6_Kernel122_Valid_Out & channel7_Kernel122_Valid_Out & channel8_Kernel122_Valid_Out & channel9_Kernel122_Valid_Out & channel10_Kernel122_Valid_Out & channel11_Kernel122_Valid_Out & channel12_Kernel122_Valid_Out & channel13_Kernel122_Valid_Out & channel14_Kernel122_Valid_Out & channel15_Kernel122_Valid_Out & channel16_Kernel122_Valid_Out & channel17_Kernel122_Valid_Out & channel18_Kernel122_Valid_Out & channel19_Kernel122_Valid_Out & channel20_Kernel122_Valid_Out & channel21_Kernel122_Valid_Out & channel22_Kernel122_Valid_Out & channel23_Kernel122_Valid_Out & channel24_Kernel122_Valid_Out & channel25_Kernel122_Valid_Out & channel26_Kernel122_Valid_Out & channel27_Kernel122_Valid_Out & channel28_Kernel122_Valid_Out & channel29_Kernel122_Valid_Out & channel30_Kernel122_Valid_Out & channel31_Kernel122_Valid_Out & channel32_Kernel122_Valid_Out & channel33_Kernel122_Valid_Out & channel34_Kernel122_Valid_Out & channel35_Kernel122_Valid_Out & channel36_Kernel122_Valid_Out & channel37_Kernel122_Valid_Out & channel38_Kernel122_Valid_Out & channel39_Kernel122_Valid_Out & channel40_Kernel122_Valid_Out & channel41_Kernel122_Valid_Out & channel42_Kernel122_Valid_Out & channel43_Kernel122_Valid_Out & channel44_Kernel122_Valid_Out & channel45_Kernel122_Valid_Out & channel46_Kernel122_Valid_Out & channel47_Kernel122_Valid_Out & channel48_Kernel122_Valid_Out & channel49_Kernel122_Valid_Out & channel50_Kernel122_Valid_Out & channel51_Kernel122_Valid_Out & channel52_Kernel122_Valid_Out & channel53_Kernel122_Valid_Out & channel54_Kernel122_Valid_Out & channel55_Kernel122_Valid_Out & channel56_Kernel122_Valid_Out & channel57_Kernel122_Valid_Out & channel58_Kernel122_Valid_Out & channel59_Kernel122_Valid_Out & channel60_Kernel122_Valid_Out & channel61_Kernel122_Valid_Out & channel62_Kernel122_Valid_Out & channel63_Kernel122_Valid_Out & channel64_Kernel122_Valid_Out;

	wire channel1_Kernel123_Valid_Out, channel2_Kernel123_Valid_Out, channel3_Kernel123_Valid_Out, channel4_Kernel123_Valid_Out, channel5_Kernel123_Valid_Out, channel6_Kernel123_Valid_Out, channel7_Kernel123_Valid_Out, channel8_Kernel123_Valid_Out, channel9_Kernel123_Valid_Out, channel10_Kernel123_Valid_Out, channel11_Kernel123_Valid_Out, channel12_Kernel123_Valid_Out, channel13_Kernel123_Valid_Out, channel14_Kernel123_Valid_Out, channel15_Kernel123_Valid_Out, channel16_Kernel123_Valid_Out, channel17_Kernel123_Valid_Out, channel18_Kernel123_Valid_Out, channel19_Kernel123_Valid_Out, channel20_Kernel123_Valid_Out, channel21_Kernel123_Valid_Out, channel22_Kernel123_Valid_Out, channel23_Kernel123_Valid_Out, channel24_Kernel123_Valid_Out, channel25_Kernel123_Valid_Out, channel26_Kernel123_Valid_Out, channel27_Kernel123_Valid_Out, channel28_Kernel123_Valid_Out, channel29_Kernel123_Valid_Out, channel30_Kernel123_Valid_Out, channel31_Kernel123_Valid_Out, channel32_Kernel123_Valid_Out, channel33_Kernel123_Valid_Out, channel34_Kernel123_Valid_Out, channel35_Kernel123_Valid_Out, channel36_Kernel123_Valid_Out, channel37_Kernel123_Valid_Out, channel38_Kernel123_Valid_Out, channel39_Kernel123_Valid_Out, channel40_Kernel123_Valid_Out, channel41_Kernel123_Valid_Out, channel42_Kernel123_Valid_Out, channel43_Kernel123_Valid_Out, channel44_Kernel123_Valid_Out, channel45_Kernel123_Valid_Out, channel46_Kernel123_Valid_Out, channel47_Kernel123_Valid_Out, channel48_Kernel123_Valid_Out, channel49_Kernel123_Valid_Out, channel50_Kernel123_Valid_Out, channel51_Kernel123_Valid_Out, channel52_Kernel123_Valid_Out, channel53_Kernel123_Valid_Out, channel54_Kernel123_Valid_Out, channel55_Kernel123_Valid_Out, channel56_Kernel123_Valid_Out, channel57_Kernel123_Valid_Out, channel58_Kernel123_Valid_Out, channel59_Kernel123_Valid_Out, channel60_Kernel123_Valid_Out, channel61_Kernel123_Valid_Out, channel62_Kernel123_Valid_Out, channel63_Kernel123_Valid_Out, channel64_Kernel123_Valid_Out;

	assign add_kernel123=channel1_Kernel123_Valid_Out & channel2_Kernel123_Valid_Out & channel3_Kernel123_Valid_Out & channel4_Kernel123_Valid_Out & channel5_Kernel123_Valid_Out & channel6_Kernel123_Valid_Out & channel7_Kernel123_Valid_Out & channel8_Kernel123_Valid_Out & channel9_Kernel123_Valid_Out & channel10_Kernel123_Valid_Out & channel11_Kernel123_Valid_Out & channel12_Kernel123_Valid_Out & channel13_Kernel123_Valid_Out & channel14_Kernel123_Valid_Out & channel15_Kernel123_Valid_Out & channel16_Kernel123_Valid_Out & channel17_Kernel123_Valid_Out & channel18_Kernel123_Valid_Out & channel19_Kernel123_Valid_Out & channel20_Kernel123_Valid_Out & channel21_Kernel123_Valid_Out & channel22_Kernel123_Valid_Out & channel23_Kernel123_Valid_Out & channel24_Kernel123_Valid_Out & channel25_Kernel123_Valid_Out & channel26_Kernel123_Valid_Out & channel27_Kernel123_Valid_Out & channel28_Kernel123_Valid_Out & channel29_Kernel123_Valid_Out & channel30_Kernel123_Valid_Out & channel31_Kernel123_Valid_Out & channel32_Kernel123_Valid_Out & channel33_Kernel123_Valid_Out & channel34_Kernel123_Valid_Out & channel35_Kernel123_Valid_Out & channel36_Kernel123_Valid_Out & channel37_Kernel123_Valid_Out & channel38_Kernel123_Valid_Out & channel39_Kernel123_Valid_Out & channel40_Kernel123_Valid_Out & channel41_Kernel123_Valid_Out & channel42_Kernel123_Valid_Out & channel43_Kernel123_Valid_Out & channel44_Kernel123_Valid_Out & channel45_Kernel123_Valid_Out & channel46_Kernel123_Valid_Out & channel47_Kernel123_Valid_Out & channel48_Kernel123_Valid_Out & channel49_Kernel123_Valid_Out & channel50_Kernel123_Valid_Out & channel51_Kernel123_Valid_Out & channel52_Kernel123_Valid_Out & channel53_Kernel123_Valid_Out & channel54_Kernel123_Valid_Out & channel55_Kernel123_Valid_Out & channel56_Kernel123_Valid_Out & channel57_Kernel123_Valid_Out & channel58_Kernel123_Valid_Out & channel59_Kernel123_Valid_Out & channel60_Kernel123_Valid_Out & channel61_Kernel123_Valid_Out & channel62_Kernel123_Valid_Out & channel63_Kernel123_Valid_Out & channel64_Kernel123_Valid_Out;

	wire channel1_Kernel124_Valid_Out, channel2_Kernel124_Valid_Out, channel3_Kernel124_Valid_Out, channel4_Kernel124_Valid_Out, channel5_Kernel124_Valid_Out, channel6_Kernel124_Valid_Out, channel7_Kernel124_Valid_Out, channel8_Kernel124_Valid_Out, channel9_Kernel124_Valid_Out, channel10_Kernel124_Valid_Out, channel11_Kernel124_Valid_Out, channel12_Kernel124_Valid_Out, channel13_Kernel124_Valid_Out, channel14_Kernel124_Valid_Out, channel15_Kernel124_Valid_Out, channel16_Kernel124_Valid_Out, channel17_Kernel124_Valid_Out, channel18_Kernel124_Valid_Out, channel19_Kernel124_Valid_Out, channel20_Kernel124_Valid_Out, channel21_Kernel124_Valid_Out, channel22_Kernel124_Valid_Out, channel23_Kernel124_Valid_Out, channel24_Kernel124_Valid_Out, channel25_Kernel124_Valid_Out, channel26_Kernel124_Valid_Out, channel27_Kernel124_Valid_Out, channel28_Kernel124_Valid_Out, channel29_Kernel124_Valid_Out, channel30_Kernel124_Valid_Out, channel31_Kernel124_Valid_Out, channel32_Kernel124_Valid_Out, channel33_Kernel124_Valid_Out, channel34_Kernel124_Valid_Out, channel35_Kernel124_Valid_Out, channel36_Kernel124_Valid_Out, channel37_Kernel124_Valid_Out, channel38_Kernel124_Valid_Out, channel39_Kernel124_Valid_Out, channel40_Kernel124_Valid_Out, channel41_Kernel124_Valid_Out, channel42_Kernel124_Valid_Out, channel43_Kernel124_Valid_Out, channel44_Kernel124_Valid_Out, channel45_Kernel124_Valid_Out, channel46_Kernel124_Valid_Out, channel47_Kernel124_Valid_Out, channel48_Kernel124_Valid_Out, channel49_Kernel124_Valid_Out, channel50_Kernel124_Valid_Out, channel51_Kernel124_Valid_Out, channel52_Kernel124_Valid_Out, channel53_Kernel124_Valid_Out, channel54_Kernel124_Valid_Out, channel55_Kernel124_Valid_Out, channel56_Kernel124_Valid_Out, channel57_Kernel124_Valid_Out, channel58_Kernel124_Valid_Out, channel59_Kernel124_Valid_Out, channel60_Kernel124_Valid_Out, channel61_Kernel124_Valid_Out, channel62_Kernel124_Valid_Out, channel63_Kernel124_Valid_Out, channel64_Kernel124_Valid_Out;

	assign add_kernel124=channel1_Kernel124_Valid_Out & channel2_Kernel124_Valid_Out & channel3_Kernel124_Valid_Out & channel4_Kernel124_Valid_Out & channel5_Kernel124_Valid_Out & channel6_Kernel124_Valid_Out & channel7_Kernel124_Valid_Out & channel8_Kernel124_Valid_Out & channel9_Kernel124_Valid_Out & channel10_Kernel124_Valid_Out & channel11_Kernel124_Valid_Out & channel12_Kernel124_Valid_Out & channel13_Kernel124_Valid_Out & channel14_Kernel124_Valid_Out & channel15_Kernel124_Valid_Out & channel16_Kernel124_Valid_Out & channel17_Kernel124_Valid_Out & channel18_Kernel124_Valid_Out & channel19_Kernel124_Valid_Out & channel20_Kernel124_Valid_Out & channel21_Kernel124_Valid_Out & channel22_Kernel124_Valid_Out & channel23_Kernel124_Valid_Out & channel24_Kernel124_Valid_Out & channel25_Kernel124_Valid_Out & channel26_Kernel124_Valid_Out & channel27_Kernel124_Valid_Out & channel28_Kernel124_Valid_Out & channel29_Kernel124_Valid_Out & channel30_Kernel124_Valid_Out & channel31_Kernel124_Valid_Out & channel32_Kernel124_Valid_Out & channel33_Kernel124_Valid_Out & channel34_Kernel124_Valid_Out & channel35_Kernel124_Valid_Out & channel36_Kernel124_Valid_Out & channel37_Kernel124_Valid_Out & channel38_Kernel124_Valid_Out & channel39_Kernel124_Valid_Out & channel40_Kernel124_Valid_Out & channel41_Kernel124_Valid_Out & channel42_Kernel124_Valid_Out & channel43_Kernel124_Valid_Out & channel44_Kernel124_Valid_Out & channel45_Kernel124_Valid_Out & channel46_Kernel124_Valid_Out & channel47_Kernel124_Valid_Out & channel48_Kernel124_Valid_Out & channel49_Kernel124_Valid_Out & channel50_Kernel124_Valid_Out & channel51_Kernel124_Valid_Out & channel52_Kernel124_Valid_Out & channel53_Kernel124_Valid_Out & channel54_Kernel124_Valid_Out & channel55_Kernel124_Valid_Out & channel56_Kernel124_Valid_Out & channel57_Kernel124_Valid_Out & channel58_Kernel124_Valid_Out & channel59_Kernel124_Valid_Out & channel60_Kernel124_Valid_Out & channel61_Kernel124_Valid_Out & channel62_Kernel124_Valid_Out & channel63_Kernel124_Valid_Out & channel64_Kernel124_Valid_Out;

	wire channel1_Kernel125_Valid_Out, channel2_Kernel125_Valid_Out, channel3_Kernel125_Valid_Out, channel4_Kernel125_Valid_Out, channel5_Kernel125_Valid_Out, channel6_Kernel125_Valid_Out, channel7_Kernel125_Valid_Out, channel8_Kernel125_Valid_Out, channel9_Kernel125_Valid_Out, channel10_Kernel125_Valid_Out, channel11_Kernel125_Valid_Out, channel12_Kernel125_Valid_Out, channel13_Kernel125_Valid_Out, channel14_Kernel125_Valid_Out, channel15_Kernel125_Valid_Out, channel16_Kernel125_Valid_Out, channel17_Kernel125_Valid_Out, channel18_Kernel125_Valid_Out, channel19_Kernel125_Valid_Out, channel20_Kernel125_Valid_Out, channel21_Kernel125_Valid_Out, channel22_Kernel125_Valid_Out, channel23_Kernel125_Valid_Out, channel24_Kernel125_Valid_Out, channel25_Kernel125_Valid_Out, channel26_Kernel125_Valid_Out, channel27_Kernel125_Valid_Out, channel28_Kernel125_Valid_Out, channel29_Kernel125_Valid_Out, channel30_Kernel125_Valid_Out, channel31_Kernel125_Valid_Out, channel32_Kernel125_Valid_Out, channel33_Kernel125_Valid_Out, channel34_Kernel125_Valid_Out, channel35_Kernel125_Valid_Out, channel36_Kernel125_Valid_Out, channel37_Kernel125_Valid_Out, channel38_Kernel125_Valid_Out, channel39_Kernel125_Valid_Out, channel40_Kernel125_Valid_Out, channel41_Kernel125_Valid_Out, channel42_Kernel125_Valid_Out, channel43_Kernel125_Valid_Out, channel44_Kernel125_Valid_Out, channel45_Kernel125_Valid_Out, channel46_Kernel125_Valid_Out, channel47_Kernel125_Valid_Out, channel48_Kernel125_Valid_Out, channel49_Kernel125_Valid_Out, channel50_Kernel125_Valid_Out, channel51_Kernel125_Valid_Out, channel52_Kernel125_Valid_Out, channel53_Kernel125_Valid_Out, channel54_Kernel125_Valid_Out, channel55_Kernel125_Valid_Out, channel56_Kernel125_Valid_Out, channel57_Kernel125_Valid_Out, channel58_Kernel125_Valid_Out, channel59_Kernel125_Valid_Out, channel60_Kernel125_Valid_Out, channel61_Kernel125_Valid_Out, channel62_Kernel125_Valid_Out, channel63_Kernel125_Valid_Out, channel64_Kernel125_Valid_Out;

	assign add_kernel125=channel1_Kernel125_Valid_Out & channel2_Kernel125_Valid_Out & channel3_Kernel125_Valid_Out & channel4_Kernel125_Valid_Out & channel5_Kernel125_Valid_Out & channel6_Kernel125_Valid_Out & channel7_Kernel125_Valid_Out & channel8_Kernel125_Valid_Out & channel9_Kernel125_Valid_Out & channel10_Kernel125_Valid_Out & channel11_Kernel125_Valid_Out & channel12_Kernel125_Valid_Out & channel13_Kernel125_Valid_Out & channel14_Kernel125_Valid_Out & channel15_Kernel125_Valid_Out & channel16_Kernel125_Valid_Out & channel17_Kernel125_Valid_Out & channel18_Kernel125_Valid_Out & channel19_Kernel125_Valid_Out & channel20_Kernel125_Valid_Out & channel21_Kernel125_Valid_Out & channel22_Kernel125_Valid_Out & channel23_Kernel125_Valid_Out & channel24_Kernel125_Valid_Out & channel25_Kernel125_Valid_Out & channel26_Kernel125_Valid_Out & channel27_Kernel125_Valid_Out & channel28_Kernel125_Valid_Out & channel29_Kernel125_Valid_Out & channel30_Kernel125_Valid_Out & channel31_Kernel125_Valid_Out & channel32_Kernel125_Valid_Out & channel33_Kernel125_Valid_Out & channel34_Kernel125_Valid_Out & channel35_Kernel125_Valid_Out & channel36_Kernel125_Valid_Out & channel37_Kernel125_Valid_Out & channel38_Kernel125_Valid_Out & channel39_Kernel125_Valid_Out & channel40_Kernel125_Valid_Out & channel41_Kernel125_Valid_Out & channel42_Kernel125_Valid_Out & channel43_Kernel125_Valid_Out & channel44_Kernel125_Valid_Out & channel45_Kernel125_Valid_Out & channel46_Kernel125_Valid_Out & channel47_Kernel125_Valid_Out & channel48_Kernel125_Valid_Out & channel49_Kernel125_Valid_Out & channel50_Kernel125_Valid_Out & channel51_Kernel125_Valid_Out & channel52_Kernel125_Valid_Out & channel53_Kernel125_Valid_Out & channel54_Kernel125_Valid_Out & channel55_Kernel125_Valid_Out & channel56_Kernel125_Valid_Out & channel57_Kernel125_Valid_Out & channel58_Kernel125_Valid_Out & channel59_Kernel125_Valid_Out & channel60_Kernel125_Valid_Out & channel61_Kernel125_Valid_Out & channel62_Kernel125_Valid_Out & channel63_Kernel125_Valid_Out & channel64_Kernel125_Valid_Out;

	wire channel1_Kernel126_Valid_Out, channel2_Kernel126_Valid_Out, channel3_Kernel126_Valid_Out, channel4_Kernel126_Valid_Out, channel5_Kernel126_Valid_Out, channel6_Kernel126_Valid_Out, channel7_Kernel126_Valid_Out, channel8_Kernel126_Valid_Out, channel9_Kernel126_Valid_Out, channel10_Kernel126_Valid_Out, channel11_Kernel126_Valid_Out, channel12_Kernel126_Valid_Out, channel13_Kernel126_Valid_Out, channel14_Kernel126_Valid_Out, channel15_Kernel126_Valid_Out, channel16_Kernel126_Valid_Out, channel17_Kernel126_Valid_Out, channel18_Kernel126_Valid_Out, channel19_Kernel126_Valid_Out, channel20_Kernel126_Valid_Out, channel21_Kernel126_Valid_Out, channel22_Kernel126_Valid_Out, channel23_Kernel126_Valid_Out, channel24_Kernel126_Valid_Out, channel25_Kernel126_Valid_Out, channel26_Kernel126_Valid_Out, channel27_Kernel126_Valid_Out, channel28_Kernel126_Valid_Out, channel29_Kernel126_Valid_Out, channel30_Kernel126_Valid_Out, channel31_Kernel126_Valid_Out, channel32_Kernel126_Valid_Out, channel33_Kernel126_Valid_Out, channel34_Kernel126_Valid_Out, channel35_Kernel126_Valid_Out, channel36_Kernel126_Valid_Out, channel37_Kernel126_Valid_Out, channel38_Kernel126_Valid_Out, channel39_Kernel126_Valid_Out, channel40_Kernel126_Valid_Out, channel41_Kernel126_Valid_Out, channel42_Kernel126_Valid_Out, channel43_Kernel126_Valid_Out, channel44_Kernel126_Valid_Out, channel45_Kernel126_Valid_Out, channel46_Kernel126_Valid_Out, channel47_Kernel126_Valid_Out, channel48_Kernel126_Valid_Out, channel49_Kernel126_Valid_Out, channel50_Kernel126_Valid_Out, channel51_Kernel126_Valid_Out, channel52_Kernel126_Valid_Out, channel53_Kernel126_Valid_Out, channel54_Kernel126_Valid_Out, channel55_Kernel126_Valid_Out, channel56_Kernel126_Valid_Out, channel57_Kernel126_Valid_Out, channel58_Kernel126_Valid_Out, channel59_Kernel126_Valid_Out, channel60_Kernel126_Valid_Out, channel61_Kernel126_Valid_Out, channel62_Kernel126_Valid_Out, channel63_Kernel126_Valid_Out, channel64_Kernel126_Valid_Out;

	assign add_kernel126=channel1_Kernel126_Valid_Out & channel2_Kernel126_Valid_Out & channel3_Kernel126_Valid_Out & channel4_Kernel126_Valid_Out & channel5_Kernel126_Valid_Out & channel6_Kernel126_Valid_Out & channel7_Kernel126_Valid_Out & channel8_Kernel126_Valid_Out & channel9_Kernel126_Valid_Out & channel10_Kernel126_Valid_Out & channel11_Kernel126_Valid_Out & channel12_Kernel126_Valid_Out & channel13_Kernel126_Valid_Out & channel14_Kernel126_Valid_Out & channel15_Kernel126_Valid_Out & channel16_Kernel126_Valid_Out & channel17_Kernel126_Valid_Out & channel18_Kernel126_Valid_Out & channel19_Kernel126_Valid_Out & channel20_Kernel126_Valid_Out & channel21_Kernel126_Valid_Out & channel22_Kernel126_Valid_Out & channel23_Kernel126_Valid_Out & channel24_Kernel126_Valid_Out & channel25_Kernel126_Valid_Out & channel26_Kernel126_Valid_Out & channel27_Kernel126_Valid_Out & channel28_Kernel126_Valid_Out & channel29_Kernel126_Valid_Out & channel30_Kernel126_Valid_Out & channel31_Kernel126_Valid_Out & channel32_Kernel126_Valid_Out & channel33_Kernel126_Valid_Out & channel34_Kernel126_Valid_Out & channel35_Kernel126_Valid_Out & channel36_Kernel126_Valid_Out & channel37_Kernel126_Valid_Out & channel38_Kernel126_Valid_Out & channel39_Kernel126_Valid_Out & channel40_Kernel126_Valid_Out & channel41_Kernel126_Valid_Out & channel42_Kernel126_Valid_Out & channel43_Kernel126_Valid_Out & channel44_Kernel126_Valid_Out & channel45_Kernel126_Valid_Out & channel46_Kernel126_Valid_Out & channel47_Kernel126_Valid_Out & channel48_Kernel126_Valid_Out & channel49_Kernel126_Valid_Out & channel50_Kernel126_Valid_Out & channel51_Kernel126_Valid_Out & channel52_Kernel126_Valid_Out & channel53_Kernel126_Valid_Out & channel54_Kernel126_Valid_Out & channel55_Kernel126_Valid_Out & channel56_Kernel126_Valid_Out & channel57_Kernel126_Valid_Out & channel58_Kernel126_Valid_Out & channel59_Kernel126_Valid_Out & channel60_Kernel126_Valid_Out & channel61_Kernel126_Valid_Out & channel62_Kernel126_Valid_Out & channel63_Kernel126_Valid_Out & channel64_Kernel126_Valid_Out;

	wire channel1_Kernel127_Valid_Out, channel2_Kernel127_Valid_Out, channel3_Kernel127_Valid_Out, channel4_Kernel127_Valid_Out, channel5_Kernel127_Valid_Out, channel6_Kernel127_Valid_Out, channel7_Kernel127_Valid_Out, channel8_Kernel127_Valid_Out, channel9_Kernel127_Valid_Out, channel10_Kernel127_Valid_Out, channel11_Kernel127_Valid_Out, channel12_Kernel127_Valid_Out, channel13_Kernel127_Valid_Out, channel14_Kernel127_Valid_Out, channel15_Kernel127_Valid_Out, channel16_Kernel127_Valid_Out, channel17_Kernel127_Valid_Out, channel18_Kernel127_Valid_Out, channel19_Kernel127_Valid_Out, channel20_Kernel127_Valid_Out, channel21_Kernel127_Valid_Out, channel22_Kernel127_Valid_Out, channel23_Kernel127_Valid_Out, channel24_Kernel127_Valid_Out, channel25_Kernel127_Valid_Out, channel26_Kernel127_Valid_Out, channel27_Kernel127_Valid_Out, channel28_Kernel127_Valid_Out, channel29_Kernel127_Valid_Out, channel30_Kernel127_Valid_Out, channel31_Kernel127_Valid_Out, channel32_Kernel127_Valid_Out, channel33_Kernel127_Valid_Out, channel34_Kernel127_Valid_Out, channel35_Kernel127_Valid_Out, channel36_Kernel127_Valid_Out, channel37_Kernel127_Valid_Out, channel38_Kernel127_Valid_Out, channel39_Kernel127_Valid_Out, channel40_Kernel127_Valid_Out, channel41_Kernel127_Valid_Out, channel42_Kernel127_Valid_Out, channel43_Kernel127_Valid_Out, channel44_Kernel127_Valid_Out, channel45_Kernel127_Valid_Out, channel46_Kernel127_Valid_Out, channel47_Kernel127_Valid_Out, channel48_Kernel127_Valid_Out, channel49_Kernel127_Valid_Out, channel50_Kernel127_Valid_Out, channel51_Kernel127_Valid_Out, channel52_Kernel127_Valid_Out, channel53_Kernel127_Valid_Out, channel54_Kernel127_Valid_Out, channel55_Kernel127_Valid_Out, channel56_Kernel127_Valid_Out, channel57_Kernel127_Valid_Out, channel58_Kernel127_Valid_Out, channel59_Kernel127_Valid_Out, channel60_Kernel127_Valid_Out, channel61_Kernel127_Valid_Out, channel62_Kernel127_Valid_Out, channel63_Kernel127_Valid_Out, channel64_Kernel127_Valid_Out;

	assign add_kernel127=channel1_Kernel127_Valid_Out & channel2_Kernel127_Valid_Out & channel3_Kernel127_Valid_Out & channel4_Kernel127_Valid_Out & channel5_Kernel127_Valid_Out & channel6_Kernel127_Valid_Out & channel7_Kernel127_Valid_Out & channel8_Kernel127_Valid_Out & channel9_Kernel127_Valid_Out & channel10_Kernel127_Valid_Out & channel11_Kernel127_Valid_Out & channel12_Kernel127_Valid_Out & channel13_Kernel127_Valid_Out & channel14_Kernel127_Valid_Out & channel15_Kernel127_Valid_Out & channel16_Kernel127_Valid_Out & channel17_Kernel127_Valid_Out & channel18_Kernel127_Valid_Out & channel19_Kernel127_Valid_Out & channel20_Kernel127_Valid_Out & channel21_Kernel127_Valid_Out & channel22_Kernel127_Valid_Out & channel23_Kernel127_Valid_Out & channel24_Kernel127_Valid_Out & channel25_Kernel127_Valid_Out & channel26_Kernel127_Valid_Out & channel27_Kernel127_Valid_Out & channel28_Kernel127_Valid_Out & channel29_Kernel127_Valid_Out & channel30_Kernel127_Valid_Out & channel31_Kernel127_Valid_Out & channel32_Kernel127_Valid_Out & channel33_Kernel127_Valid_Out & channel34_Kernel127_Valid_Out & channel35_Kernel127_Valid_Out & channel36_Kernel127_Valid_Out & channel37_Kernel127_Valid_Out & channel38_Kernel127_Valid_Out & channel39_Kernel127_Valid_Out & channel40_Kernel127_Valid_Out & channel41_Kernel127_Valid_Out & channel42_Kernel127_Valid_Out & channel43_Kernel127_Valid_Out & channel44_Kernel127_Valid_Out & channel45_Kernel127_Valid_Out & channel46_Kernel127_Valid_Out & channel47_Kernel127_Valid_Out & channel48_Kernel127_Valid_Out & channel49_Kernel127_Valid_Out & channel50_Kernel127_Valid_Out & channel51_Kernel127_Valid_Out & channel52_Kernel127_Valid_Out & channel53_Kernel127_Valid_Out & channel54_Kernel127_Valid_Out & channel55_Kernel127_Valid_Out & channel56_Kernel127_Valid_Out & channel57_Kernel127_Valid_Out & channel58_Kernel127_Valid_Out & channel59_Kernel127_Valid_Out & channel60_Kernel127_Valid_Out & channel61_Kernel127_Valid_Out & channel62_Kernel127_Valid_Out & channel63_Kernel127_Valid_Out & channel64_Kernel127_Valid_Out;

	wire channel1_Kernel128_Valid_Out, channel2_Kernel128_Valid_Out, channel3_Kernel128_Valid_Out, channel4_Kernel128_Valid_Out, channel5_Kernel128_Valid_Out, channel6_Kernel128_Valid_Out, channel7_Kernel128_Valid_Out, channel8_Kernel128_Valid_Out, channel9_Kernel128_Valid_Out, channel10_Kernel128_Valid_Out, channel11_Kernel128_Valid_Out, channel12_Kernel128_Valid_Out, channel13_Kernel128_Valid_Out, channel14_Kernel128_Valid_Out, channel15_Kernel128_Valid_Out, channel16_Kernel128_Valid_Out, channel17_Kernel128_Valid_Out, channel18_Kernel128_Valid_Out, channel19_Kernel128_Valid_Out, channel20_Kernel128_Valid_Out, channel21_Kernel128_Valid_Out, channel22_Kernel128_Valid_Out, channel23_Kernel128_Valid_Out, channel24_Kernel128_Valid_Out, channel25_Kernel128_Valid_Out, channel26_Kernel128_Valid_Out, channel27_Kernel128_Valid_Out, channel28_Kernel128_Valid_Out, channel29_Kernel128_Valid_Out, channel30_Kernel128_Valid_Out, channel31_Kernel128_Valid_Out, channel32_Kernel128_Valid_Out, channel33_Kernel128_Valid_Out, channel34_Kernel128_Valid_Out, channel35_Kernel128_Valid_Out, channel36_Kernel128_Valid_Out, channel37_Kernel128_Valid_Out, channel38_Kernel128_Valid_Out, channel39_Kernel128_Valid_Out, channel40_Kernel128_Valid_Out, channel41_Kernel128_Valid_Out, channel42_Kernel128_Valid_Out, channel43_Kernel128_Valid_Out, channel44_Kernel128_Valid_Out, channel45_Kernel128_Valid_Out, channel46_Kernel128_Valid_Out, channel47_Kernel128_Valid_Out, channel48_Kernel128_Valid_Out, channel49_Kernel128_Valid_Out, channel50_Kernel128_Valid_Out, channel51_Kernel128_Valid_Out, channel52_Kernel128_Valid_Out, channel53_Kernel128_Valid_Out, channel54_Kernel128_Valid_Out, channel55_Kernel128_Valid_Out, channel56_Kernel128_Valid_Out, channel57_Kernel128_Valid_Out, channel58_Kernel128_Valid_Out, channel59_Kernel128_Valid_Out, channel60_Kernel128_Valid_Out, channel61_Kernel128_Valid_Out, channel62_Kernel128_Valid_Out, channel63_Kernel128_Valid_Out, channel64_Kernel128_Valid_Out;

	assign add_kernel128=channel1_Kernel128_Valid_Out & channel2_Kernel128_Valid_Out & channel3_Kernel128_Valid_Out & channel4_Kernel128_Valid_Out & channel5_Kernel128_Valid_Out & channel6_Kernel128_Valid_Out & channel7_Kernel128_Valid_Out & channel8_Kernel128_Valid_Out & channel9_Kernel128_Valid_Out & channel10_Kernel128_Valid_Out & channel11_Kernel128_Valid_Out & channel12_Kernel128_Valid_Out & channel13_Kernel128_Valid_Out & channel14_Kernel128_Valid_Out & channel15_Kernel128_Valid_Out & channel16_Kernel128_Valid_Out & channel17_Kernel128_Valid_Out & channel18_Kernel128_Valid_Out & channel19_Kernel128_Valid_Out & channel20_Kernel128_Valid_Out & channel21_Kernel128_Valid_Out & channel22_Kernel128_Valid_Out & channel23_Kernel128_Valid_Out & channel24_Kernel128_Valid_Out & channel25_Kernel128_Valid_Out & channel26_Kernel128_Valid_Out & channel27_Kernel128_Valid_Out & channel28_Kernel128_Valid_Out & channel29_Kernel128_Valid_Out & channel30_Kernel128_Valid_Out & channel31_Kernel128_Valid_Out & channel32_Kernel128_Valid_Out & channel33_Kernel128_Valid_Out & channel34_Kernel128_Valid_Out & channel35_Kernel128_Valid_Out & channel36_Kernel128_Valid_Out & channel37_Kernel128_Valid_Out & channel38_Kernel128_Valid_Out & channel39_Kernel128_Valid_Out & channel40_Kernel128_Valid_Out & channel41_Kernel128_Valid_Out & channel42_Kernel128_Valid_Out & channel43_Kernel128_Valid_Out & channel44_Kernel128_Valid_Out & channel45_Kernel128_Valid_Out & channel46_Kernel128_Valid_Out & channel47_Kernel128_Valid_Out & channel48_Kernel128_Valid_Out & channel49_Kernel128_Valid_Out & channel50_Kernel128_Valid_Out & channel51_Kernel128_Valid_Out & channel52_Kernel128_Valid_Out & channel53_Kernel128_Valid_Out & channel54_Kernel128_Valid_Out & channel55_Kernel128_Valid_Out & channel56_Kernel128_Valid_Out & channel57_Kernel128_Valid_Out & channel58_Kernel128_Valid_Out & channel59_Kernel128_Valid_Out & channel60_Kernel128_Valid_Out & channel61_Kernel128_Valid_Out & channel62_Kernel128_Valid_Out & channel63_Kernel128_Valid_Out & channel64_Kernel128_Valid_Out;


	wire [31:0] bn1_Data_Out, bn2_Data_Out, bn3_Data_Out, bn4_Data_Out, bn5_Data_Out, bn6_Data_Out, bn7_Data_Out, bn8_Data_Out, bn9_Data_Out, bn10_Data_Out, bn11_Data_Out, bn12_Data_Out, bn13_Data_Out, bn14_Data_Out, bn15_Data_Out, bn16_Data_Out, bn17_Data_Out, bn18_Data_Out, bn19_Data_Out, bn20_Data_Out, bn21_Data_Out, bn22_Data_Out, bn23_Data_Out, bn24_Data_Out, bn25_Data_Out, bn26_Data_Out, bn27_Data_Out, bn28_Data_Out, bn29_Data_Out, bn30_Data_Out, bn31_Data_Out, bn32_Data_Out, bn33_Data_Out, bn34_Data_Out, bn35_Data_Out, bn36_Data_Out, bn37_Data_Out, bn38_Data_Out, bn39_Data_Out, bn40_Data_Out, bn41_Data_Out, bn42_Data_Out, bn43_Data_Out, bn44_Data_Out, bn45_Data_Out, bn46_Data_Out, bn47_Data_Out, bn48_Data_Out, bn49_Data_Out, bn50_Data_Out, bn51_Data_Out, bn52_Data_Out, bn53_Data_Out, bn54_Data_Out, bn55_Data_Out, bn56_Data_Out, bn57_Data_Out, bn58_Data_Out, bn59_Data_Out, bn60_Data_Out, bn61_Data_Out, bn62_Data_Out, bn63_Data_Out, bn64_Data_Out, bn65_Data_Out, bn66_Data_Out, bn67_Data_Out, bn68_Data_Out, bn69_Data_Out, bn70_Data_Out, bn71_Data_Out, bn72_Data_Out, bn73_Data_Out, bn74_Data_Out, bn75_Data_Out, bn76_Data_Out, bn77_Data_Out, bn78_Data_Out, bn79_Data_Out, bn80_Data_Out, bn81_Data_Out, bn82_Data_Out, bn83_Data_Out, bn84_Data_Out, bn85_Data_Out, bn86_Data_Out, bn87_Data_Out, bn88_Data_Out, bn89_Data_Out, bn90_Data_Out, bn91_Data_Out, bn92_Data_Out, bn93_Data_Out, bn94_Data_Out, bn95_Data_Out, bn96_Data_Out, bn97_Data_Out, bn98_Data_Out, bn99_Data_Out, bn100_Data_Out, bn101_Data_Out, bn102_Data_Out, bn103_Data_Out, bn104_Data_Out, bn105_Data_Out, bn106_Data_Out, bn107_Data_Out, bn108_Data_Out, bn109_Data_Out, bn110_Data_Out, bn111_Data_Out, bn112_Data_Out, bn113_Data_Out, bn114_Data_Out, bn115_Data_Out, bn116_Data_Out, bn117_Data_Out, bn118_Data_Out, bn119_Data_Out, bn120_Data_Out, bn121_Data_Out, bn122_Data_Out, bn123_Data_Out, bn124_Data_Out, bn125_Data_Out, bn126_Data_Out, bn127_Data_Out, bn128_Data_Out;

	wire bn1_Valid_Out, bn2_Valid_Out, bn3_Valid_Out, bn4_Valid_Out, bn5_Valid_Out, bn6_Valid_Out, bn7_Valid_Out, bn8_Valid_Out, bn9_Valid_Out, bn10_Valid_Out, bn11_Valid_Out, bn12_Valid_Out, bn13_Valid_Out, bn14_Valid_Out, bn15_Valid_Out, bn16_Valid_Out, bn17_Valid_Out, bn18_Valid_Out, bn19_Valid_Out, bn20_Valid_Out, bn21_Valid_Out, bn22_Valid_Out, bn23_Valid_Out, bn24_Valid_Out, bn25_Valid_Out, bn26_Valid_Out, bn27_Valid_Out, bn28_Valid_Out, bn29_Valid_Out, bn30_Valid_Out, bn31_Valid_Out, bn32_Valid_Out, bn33_Valid_Out, bn34_Valid_Out, bn35_Valid_Out, bn36_Valid_Out, bn37_Valid_Out, bn38_Valid_Out, bn39_Valid_Out, bn40_Valid_Out, bn41_Valid_Out, bn42_Valid_Out, bn43_Valid_Out, bn44_Valid_Out, bn45_Valid_Out, bn46_Valid_Out, bn47_Valid_Out, bn48_Valid_Out, bn49_Valid_Out, bn50_Valid_Out, bn51_Valid_Out, bn52_Valid_Out, bn53_Valid_Out, bn54_Valid_Out, bn55_Valid_Out, bn56_Valid_Out, bn57_Valid_Out, bn58_Valid_Out, bn59_Valid_Out, bn60_Valid_Out, bn61_Valid_Out, bn62_Valid_Out, bn63_Valid_Out, bn64_Valid_Out, bn65_Valid_Out, bn66_Valid_Out, bn67_Valid_Out, bn68_Valid_Out, bn69_Valid_Out, bn70_Valid_Out, bn71_Valid_Out, bn72_Valid_Out, bn73_Valid_Out, bn74_Valid_Out, bn75_Valid_Out, bn76_Valid_Out, bn77_Valid_Out, bn78_Valid_Out, bn79_Valid_Out, bn80_Valid_Out, bn81_Valid_Out, bn82_Valid_Out, bn83_Valid_Out, bn84_Valid_Out, bn85_Valid_Out, bn86_Valid_Out, bn87_Valid_Out, bn88_Valid_Out, bn89_Valid_Out, bn90_Valid_Out, bn91_Valid_Out, bn92_Valid_Out, bn93_Valid_Out, bn94_Valid_Out, bn95_Valid_Out, bn96_Valid_Out, bn97_Valid_Out, bn98_Valid_Out, bn99_Valid_Out, bn100_Valid_Out, bn101_Valid_Out, bn102_Valid_Out, bn103_Valid_Out, bn104_Valid_Out, bn105_Valid_Out, bn106_Valid_Out, bn107_Valid_Out, bn108_Valid_Out, bn109_Valid_Out, bn110_Valid_Out, bn111_Valid_Out, bn112_Valid_Out, bn113_Valid_Out, bn114_Valid_Out, bn115_Valid_Out, bn116_Valid_Out, bn117_Valid_Out, bn118_Valid_Out, bn119_Valid_Out, bn120_Valid_Out, bn121_Valid_Out, bn122_Valid_Out, bn123_Valid_Out, bn124_Valid_Out, bn125_Valid_Out, bn126_Valid_Out, bn127_Valid_Out, bn128_Valid_Out;

	wire rl1_Valid_Out, rl2_Valid_Out, rl3_Valid_Out, rl4_Valid_Out, rl5_Valid_Out, rl6_Valid_Out, rl7_Valid_Out, rl8_Valid_Out, rl9_Valid_Out, rl10_Valid_Out, rl11_Valid_Out, rl12_Valid_Out, rl13_Valid_Out, rl14_Valid_Out, rl15_Valid_Out, rl16_Valid_Out, rl17_Valid_Out, rl18_Valid_Out, rl19_Valid_Out, rl20_Valid_Out, rl21_Valid_Out, rl22_Valid_Out, rl23_Valid_Out, rl24_Valid_Out, rl25_Valid_Out, rl26_Valid_Out, rl27_Valid_Out, rl28_Valid_Out, rl29_Valid_Out, rl30_Valid_Out, rl31_Valid_Out, rl32_Valid_Out, rl33_Valid_Out, rl34_Valid_Out, rl35_Valid_Out, rl36_Valid_Out, rl37_Valid_Out, rl38_Valid_Out, rl39_Valid_Out, rl40_Valid_Out, rl41_Valid_Out, rl42_Valid_Out, rl43_Valid_Out, rl44_Valid_Out, rl45_Valid_Out, rl46_Valid_Out, rl47_Valid_Out, rl48_Valid_Out, rl49_Valid_Out, rl50_Valid_Out, rl51_Valid_Out, rl52_Valid_Out, rl53_Valid_Out, rl54_Valid_Out, rl55_Valid_Out, rl56_Valid_Out, rl57_Valid_Out, rl58_Valid_Out, rl59_Valid_Out, rl60_Valid_Out, rl61_Valid_Out, rl62_Valid_Out, rl63_Valid_Out, rl64_Valid_Out, rl65_Valid_Out, rl66_Valid_Out, rl67_Valid_Out, rl68_Valid_Out, rl69_Valid_Out, rl70_Valid_Out, rl71_Valid_Out, rl72_Valid_Out, rl73_Valid_Out, rl74_Valid_Out, rl75_Valid_Out, rl76_Valid_Out, rl77_Valid_Out, rl78_Valid_Out, rl79_Valid_Out, rl80_Valid_Out, rl81_Valid_Out, rl82_Valid_Out, rl83_Valid_Out, rl84_Valid_Out, rl85_Valid_Out, rl86_Valid_Out, rl87_Valid_Out, rl88_Valid_Out, rl89_Valid_Out, rl90_Valid_Out, rl91_Valid_Out, rl92_Valid_Out, rl93_Valid_Out, rl94_Valid_Out, rl95_Valid_Out, rl96_Valid_Out, rl97_Valid_Out, rl98_Valid_Out, rl99_Valid_Out, rl100_Valid_Out, rl101_Valid_Out, rl102_Valid_Out, rl103_Valid_Out, rl104_Valid_Out, rl105_Valid_Out, rl106_Valid_Out, rl107_Valid_Out, rl108_Valid_Out, rl109_Valid_Out, rl110_Valid_Out, rl111_Valid_Out, rl112_Valid_Out, rl113_Valid_Out, rl114_Valid_Out, rl115_Valid_Out, rl116_Valid_Out, rl117_Valid_Out, rl118_Valid_Out, rl119_Valid_Out, rl120_Valid_Out, rl121_Valid_Out, rl122_Valid_Out, rl123_Valid_Out, rl124_Valid_Out, rl125_Valid_Out, rl126_Valid_Out, rl127_Valid_Out, rl128_Valid_Out;

	 assign Valid_Out = rl1_Valid_Out & rl2_Valid_Out & rl3_Valid_Out & rl4_Valid_Out & rl5_Valid_Out & rl6_Valid_Out & rl7_Valid_Out & rl8_Valid_Out & rl9_Valid_Out & rl10_Valid_Out & rl11_Valid_Out & rl12_Valid_Out & rl13_Valid_Out & rl14_Valid_Out & rl15_Valid_Out & rl16_Valid_Out & rl17_Valid_Out & rl18_Valid_Out & rl19_Valid_Out & rl20_Valid_Out & rl21_Valid_Out & rl22_Valid_Out & rl23_Valid_Out & rl24_Valid_Out & rl25_Valid_Out & rl26_Valid_Out & rl27_Valid_Out & rl28_Valid_Out & rl29_Valid_Out & rl30_Valid_Out & rl31_Valid_Out & rl32_Valid_Out & rl33_Valid_Out & rl34_Valid_Out & rl35_Valid_Out & rl36_Valid_Out & rl37_Valid_Out & rl38_Valid_Out & rl39_Valid_Out & rl40_Valid_Out & rl41_Valid_Out & rl42_Valid_Out & rl43_Valid_Out & rl44_Valid_Out & rl45_Valid_Out & rl46_Valid_Out & rl47_Valid_Out & rl48_Valid_Out & rl49_Valid_Out & rl50_Valid_Out & rl51_Valid_Out & rl52_Valid_Out & rl53_Valid_Out & rl54_Valid_Out & rl55_Valid_Out & rl56_Valid_Out & rl57_Valid_Out & rl58_Valid_Out & rl59_Valid_Out & rl60_Valid_Out & rl61_Valid_Out & rl62_Valid_Out & rl63_Valid_Out & rl64_Valid_Out & rl65_Valid_Out & rl66_Valid_Out & rl67_Valid_Out & rl68_Valid_Out & rl69_Valid_Out & rl70_Valid_Out & rl71_Valid_Out & rl72_Valid_Out & rl73_Valid_Out & rl74_Valid_Out & rl75_Valid_Out & rl76_Valid_Out & rl77_Valid_Out & rl78_Valid_Out & rl79_Valid_Out & rl80_Valid_Out & rl81_Valid_Out & rl82_Valid_Out & rl83_Valid_Out & rl84_Valid_Out & rl85_Valid_Out & rl86_Valid_Out & rl87_Valid_Out & rl88_Valid_Out & rl89_Valid_Out & rl90_Valid_Out & rl91_Valid_Out & rl92_Valid_Out & rl93_Valid_Out & rl94_Valid_Out & rl95_Valid_Out & rl96_Valid_Out & rl97_Valid_Out & rl98_Valid_Out & rl99_Valid_Out & rl100_Valid_Out & rl101_Valid_Out & rl102_Valid_Out & rl103_Valid_Out & rl104_Valid_Out & rl105_Valid_Out & rl106_Valid_Out & rl107_Valid_Out & rl108_Valid_Out & rl109_Valid_Out & rl110_Valid_Out & rl111_Valid_Out & rl112_Valid_Out & rl113_Valid_Out & rl114_Valid_Out & rl115_Valid_Out & rl116_Valid_Out & rl117_Valid_Out & rl118_Valid_Out & rl119_Valid_Out & rl120_Valid_Out & rl121_Valid_Out & rl122_Valid_Out & rl123_Valid_Out & rl124_Valid_Out & rl125_Valid_Out & rl126_Valid_Out & rl127_Valid_Out & rl128_Valid_Out;
//////////KERNEL1//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111110100110101011111101000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111100110110010111011100010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110001010000110100011001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110101111100101000111000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111101100101111001100010110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111101110001011110100110111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111101100101000111001001001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111101001101100011100101101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111101100101000100011001010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111010110110000101010111010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111100110101001101110100000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111101001101100001011010100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111101100111111010000101100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111110100101101111101101011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110101010011011111110111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111011100100100001001001010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111111001001001101010100010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111101011110000101110011011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110001010100010011100000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110100111000001101001000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110101101000111100101000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111110000110110100101010100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110000100000010111011001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111110100010010100111000111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111110100010100010110010110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110001101000010010010100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110000110110100110101110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111110001000100111101100010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111110011000010000011100101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111110010001101110000011011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111100010100101011100100000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110110011101010011000010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111101101011000010000100101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b00111110001111111111111100000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111110101110110101111101100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b10111100110001000100011110011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111101010001000101101101000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b00111101000000101111001001000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b00111110011110111100011010100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111101000011010111001010011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111110111101100111100110110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111110100111111110101001000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111011100111111000101000101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b00111011111110100001100111001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111110100111110000110011100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111110010011011001101001001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111110010010001011000000011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111110110001001000010011000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111101101100111100110001100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111100111110010110010000010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111110010001111001110110011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111110001000001111110011001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b00111110000100011011011111110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111110110111110111110101011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b10111101111110001001100101110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111101110000011011100011010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111110110000011111011110100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b10111101100111101111001010001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111101100001000011011110101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111100101111001000001011110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111110010010111101000100010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b10111110000010000111111101100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111101010110001111000100111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b10111101000010101100100101011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel1_Valid_Out)
	);
	Adder_64input add_k1(
		.Data1(Data_Out_Kernel1[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel1[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel1[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel1[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel1[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel1[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel1[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel1[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel1[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel1[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel1[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel1[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel1[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel1[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel1[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel1[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel1[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel1[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel1[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel1[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel1[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel1[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel1[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel1[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel1[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel1[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel1[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel1[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel1[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel1[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel1[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel1[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel1[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel1[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel1[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel1[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel1[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel1[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel1[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel1[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel1[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel1[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel1[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel1[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel1[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel1[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel1[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel1[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel1[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel1[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel1[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel1[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel1[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel1[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel1[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel1[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel1[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel1[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel1[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel1[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel1[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel1[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel1[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel1[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel1),
		.Data_Out(add_k1_Data_Out),
		.Valid_Out(add_kernel1_Valid_Out)
	);
	Batch_Norm bn_kernel1(
		.Data_A(32'b00111110010101101101111000100000),
		.Data_B(32'b10111111011011001011011100011011),
		.Data_In(add_k1_Data_Out),
		.Valid_In(add_kernel1_Valid_Out),
		.Data_Out(bn1_Data_Out),
		.Valid_Out(bn1_Valid_Out)
	);
	Relu_Core rl_kernel1(
		.Data_In(bn1_Data_Out),
		.Valid_In(bn1_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT-1:0]),
		.Valid_Out(rl1_Valid_Out)
	);
//////////KERNEL2//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110110101011111111101110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111110111101100110000111011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110101110011011010111101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110111001111010000101001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111110000001101110110010110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111101101101100111011100001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111110000101011010010100010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111101110010011010010000010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111110101011110111001100111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111101111111100000001000101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111100000101000110101011100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110100001011010000011001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111101111000110010101011011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111100011000111111011000011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110110100110100101100000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111100111110101111011010010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111110111000010000110111010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111101001000110101100101110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111100100001000010100110100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111100100000101010100101001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110100111101100001110000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111101010101111010111110001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111110111001100110110100010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111110001010000010000001101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111101111001111101010011101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111110011101100111110110100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111110100000010111000010000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111110101100011001011100111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111110100101110111001100000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110100011001111111010110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111110000111010101010110000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111110110000010001110011101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b00111110000110011110001101011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111110010110111000010001110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111110100100000001111110010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111110010101000111010100001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b10111110101111110011101000111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111110000101110100000110101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111110010000101010111101100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b00111100001101110011010000011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b10111111001100010011000000111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b10111101101111101001000000001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b00111110000010101011010110101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b00111101010101010011100011101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b00111101100000000010111111010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b10111110100011110110111000100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b10111101111011000101111100101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b00111110001111111100011111011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b00111101100110011000000100011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111101111001111111001000100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111101011010111111000001000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b10111110001110101011100011011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111110001100000000011011100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b00111101010110101101000000111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b10111101101101101101011010001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111101110100001100110100010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b10111110010101001100000100110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b10111110101101111111101111011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111100001111001010110011101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111101110010110100010010000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b10111110011001001110101110011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111011111110000001111110111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111101111010101001100100100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111110100110110010111110100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel2_Valid_Out)
	);
	Adder_64input add_k2(
		.Data1(Data_Out_Kernel2[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel2[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel2[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel2[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel2[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel2[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel2[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel2[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel2[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel2[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel2[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel2[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel2[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel2[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel2[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel2[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel2[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel2[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel2[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel2[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel2[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel2[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel2[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel2[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel2[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel2[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel2[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel2[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel2[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel2[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel2[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel2[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel2[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel2[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel2[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel2[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel2[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel2[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel2[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel2[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel2[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel2[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel2[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel2[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel2[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel2[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel2[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel2[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel2[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel2[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel2[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel2[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel2[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel2[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel2[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel2[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel2[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel2[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel2[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel2[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel2[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel2[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel2[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel2[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel2),
		.Data_Out(add_k2_Data_Out),
		.Valid_Out(add_kernel2_Valid_Out)
	);
	Batch_Norm bn_kernel2(
		.Data_A(32'b00111110010000010111101010011111),
		.Data_B(32'b00111111001110110010110011011111),
		.Data_In(add_k2_Data_Out),
		.Valid_In(add_kernel2_Valid_Out),
		.Data_Out(bn2_Data_Out),
		.Valid_Out(bn2_Valid_Out)
	);
	Relu_Core rl_kernel2(
		.Data_In(bn2_Data_Out),
		.Valid_In(bn2_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Valid_Out(rl2_Valid_Out)
	);
//////////KERNEL3//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110101011111000111101101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111110100110110001111011011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110011001011001101100001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110011011110100011001011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111101101011001100110110000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111011011101001011011001011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111110011100101001010011100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111101111011011010100001110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111110011110100110110001001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110001101110110011100101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111100101011000001000101010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110000010010011010000100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111101101111011100000010110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111110000111100110110000101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110101110111001111101100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111110101000111111111010011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111101100101010011010011100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111110010110010100000000111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111110000000101001001011000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111100011111110100000011001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110101010000111010111100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111110000100011110111110101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111110110111011101000101011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111110001001011011011110110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111110001110011111011011011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111110011011011000001010001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111111000100100110111111011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111111000011011110000100001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111101010010011010000001110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111111000111010011110011101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111110011101110001001100011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111100001001011010110001010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111101000001101011111111110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111110111111111011000001000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111111001111111000011001100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111110011000010111001111000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111101000111110001010010110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b00111101011011111111001101110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111110010010000110111110010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111101010111011010101111011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b10111110111101101010001110010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111101001110000111000001000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b00111101011001001010101110000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b00111110000000100011100011001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b00111110011001011110101000100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b10111110100000111101010101010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b10111101110100100001010110000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b00111110101101100111010010011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b00111110000000000000011110100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b00111110000011100000010001111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111100100111010010110011110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b10111110011100010100010001110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111101101110100101111111110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b00111101101001110100111000000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b10111110000011000110100001011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b00111101110101110011000001110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b10111110000101111010111010110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b10111110101000011000100011110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111110101110111001101110000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b00111100100100100011111100010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111101011000100101110000111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111101100010011110110111010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b10111110000101100101000110101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111110100001010111000111101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel3_Valid_Out)
	);
	Adder_64input add_k3(
		.Data1(Data_Out_Kernel3[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel3[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel3[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel3[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel3[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel3[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel3[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel3[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel3[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel3[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel3[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel3[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel3[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel3[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel3[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel3[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel3[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel3[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel3[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel3[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel3[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel3[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel3[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel3[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel3[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel3[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel3[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel3[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel3[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel3[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel3[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel3[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel3[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel3[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel3[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel3[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel3[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel3[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel3[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel3[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel3[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel3[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel3[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel3[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel3[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel3[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel3[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel3[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel3[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel3[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel3[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel3[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel3[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel3[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel3[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel3[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel3[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel3[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel3[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel3[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel3[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel3[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel3[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel3[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel3),
		.Data_Out(add_k3_Data_Out),
		.Valid_Out(add_kernel3_Valid_Out)
	);
	Batch_Norm bn_kernel3(
		.Data_A(32'b00111110011010010010110101100111),
		.Data_B(32'b10111101000011010000000101001000),
		.Data_In(add_k3_Data_Out),
		.Valid_In(add_kernel3_Valid_Out),
		.Data_Out(bn3_Data_Out),
		.Valid_Out(bn3_Valid_Out)
	);
	Relu_Core rl_kernel3(
		.Data_In(bn3_Data_Out),
		.Valid_In(bn3_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(rl3_Valid_Out)
	);
//////////KERNEL4//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111110111001001000111111001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110101110000110101010001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111101111011110011010101111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111100100100001010011111000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111110000110111100100110001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111101101110100001101010101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111110100110011001110101010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111101001000100100000100100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111100101101101110000011111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111110011100011110001000110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111101100010110110011100100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111101110001000000000110111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111101110011000110011010101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111101010001011010011001100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110000110010010110011001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111110100101101110011011100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111100001011111100101010010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110100001100010110000110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110100001001110000100011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111101100001000100001110010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110101101000011010001000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111110011010101101010111110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110011001101110000100100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111110000010111001111000111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111110011100011111000110111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110101110110110011111010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111111000111011100010010011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110001111111000011101010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111101101111100101001101010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111110101001001000110100110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111110110100000000100111100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110100110111100110011000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b00111110100000110111010000001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b00111110100101111001111011010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111110110100101110110101111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111100101100000000001100010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111100110001011010110001000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111110000100101110010001011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b00111101110000101001101010010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b00111100110001111011101010010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111111001110011010100001101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111100110100101001111100001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111101010001000111110110010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111110110010100001010000001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111101100111010000100111100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111110110101100110100100000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111110011101101111110110111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111110100011101011001010100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b00111100101011100011011100101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111101100010011000010110001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111100110101110100010111011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111110000000000010000110010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b00111101111000101001001010011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111110100100011111110111100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111101101001101111101100010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111101100011110101111011011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111110010111111111100101101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111110100111111110011000000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b10111110010111000001110011011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111100101010100010001000010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b10111101000100111010111100111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111101000110101111001110110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111110111001011011000101011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b10111110000100011001101101001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel4_Valid_Out)
	);
	Adder_64input add_k4(
		.Data1(Data_Out_Kernel4[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel4[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel4[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel4[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel4[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel4[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel4[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel4[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel4[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel4[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel4[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel4[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel4[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel4[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel4[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel4[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel4[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel4[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel4[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel4[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel4[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel4[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel4[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel4[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel4[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel4[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel4[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel4[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel4[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel4[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel4[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel4[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel4[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel4[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel4[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel4[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel4[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel4[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel4[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel4[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel4[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel4[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel4[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel4[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel4[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel4[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel4[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel4[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel4[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel4[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel4[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel4[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel4[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel4[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel4[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel4[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel4[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel4[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel4[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel4[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel4[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel4[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel4[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel4[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel4),
		.Data_Out(add_k4_Data_Out),
		.Valid_Out(add_kernel4_Valid_Out)
	);
	Batch_Norm bn_kernel4(
		.Data_A(32'b00111110011101100100111011100010),
		.Data_B(32'b10111110001101011011011011100001),
		.Data_In(add_k4_Data_Out),
		.Valid_In(add_kernel4_Valid_Out),
		.Data_Out(bn4_Data_Out),
		.Valid_Out(bn4_Valid_Out)
	);
	Relu_Core rl_kernel4(
		.Data_In(bn4_Data_Out),
		.Valid_In(bn4_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(rl4_Valid_Out)
	);
//////////KERNEL5//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111110101000011001010001011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111100100101000111101010000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110110010010000111110101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110011001101000101101101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111110010111101000011000000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110010001100100111111000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111111100010010001000100011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111110110001001011100011011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111100110000010101100000100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111110101000001100101001010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111101101011001001111000000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111110110011011101010100011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111110000000010111011111000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111110000010011000001001010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110100100101100111101100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111110011101001000110101010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111111000100101100110100111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111110010010110111101101100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111110000010000110101110001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110101011110110100101111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111100110101000111011100101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111110101000100000000011011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110101110001010101100100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111110010101100111010001111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111110111111111101011010010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111101110010010110100001101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110010001001110111110000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111101000011111000100101111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111110100010100101111111101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111110110010010000000111101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111110010011111100101010111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110011111110111010001000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b00111110100011010010010110100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b00111110101000001011010111001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111111010111001100101101100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b10111110110000000010000111011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111110110000000010000001011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b00111110010010111111010100111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111101101111011010101010011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111110010000100011110111101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b10111101100100001001001000011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b10111110100100100010110010101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b00111101000110111001110111000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b00111101100101001101011101000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111110110000100100110000001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111110100000110100010010110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111110000111101011001000000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111110101011110000100010000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111111000100010110001111110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b00111101111101001111000011110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111101111110001110110010010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111110000110111101011100001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b00111111001010010010001100110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b00111110100111011100100111111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b10111100100001110100001010111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111110101101011111100010001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111111010000000001100111010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111101011111110000110001111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b10111110011011001000001110111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b00111111000111100010011001011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111101111011110100100101111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b10111110000001011100010100001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111101110110111000001110011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111110101000001101100111101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel5_Valid_Out)
	);
	Adder_64input add_k5(
		.Data1(Data_Out_Kernel5[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel5[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel5[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel5[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel5[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel5[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel5[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel5[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel5[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel5[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel5[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel5[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel5[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel5[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel5[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel5[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel5[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel5[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel5[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel5[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel5[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel5[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel5[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel5[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel5[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel5[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel5[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel5[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel5[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel5[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel5[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel5[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel5[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel5[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel5[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel5[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel5[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel5[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel5[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel5[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel5[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel5[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel5[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel5[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel5[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel5[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel5[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel5[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel5[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel5[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel5[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel5[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel5[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel5[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel5[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel5[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel5[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel5[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel5[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel5[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel5[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel5[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel5[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel5[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel5),
		.Data_Out(add_k5_Data_Out),
		.Valid_Out(add_kernel5_Valid_Out)
	);
	Batch_Norm bn_kernel5(
		.Data_A(32'b00111110001000111011101011001100),
		.Data_B(32'b10111101110101000100100010111101),
		.Data_In(add_k5_Data_Out),
		.Valid_In(add_kernel5_Valid_Out),
		.Data_Out(bn5_Data_Out),
		.Valid_Out(bn5_Valid_Out)
	);
	Relu_Core rl_kernel5(
		.Data_In(bn5_Data_Out),
		.Valid_In(bn5_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(rl5_Valid_Out)
	);
//////////KERNEL6//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111111000000000010100101000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111101100001110110010111100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110010111010011000111001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110010010000111100000101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111101011111011101111111110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111100110011110010111111101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111110100001111011011110001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111101110001001100101110101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110011100000111101001000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111110000000100110010110010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111101111110011010011000010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111110011000110010011010000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110001101101100100001011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111101101110101010010110000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110100111011100111011010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111010111001010101110110011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110100000110110100100110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111101000011111111011110101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110011011110010011010100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110101111101000100101111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110010000110001010010010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111100011001101010010101111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110110110011110100110110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111110000001001011101111010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111110100011100001011000110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110010101001100010001001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110011100011010111111111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110011000101111000000111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111101100000011100011110111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111110100010011001000111011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111101101101110101100110110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111101111001110000000001001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b00111100011110000001101111101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b00111110100011001111001000101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111111000010011010001110010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b10111100111111100100001010100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111110101100011110100011100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111100100100110000100101010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b00111101100110001101111100010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111101111011110101000010100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111111000001101000110000000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111100111111111110010010000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111101110011000000011101010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111110001000001111111011011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111101100110010111101101110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111110100001000010001011011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111110101011100101011110100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111110101110110000011000010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111101000100000100010101101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111101011001000101101101100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111101101001111011111011110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111110001000100000010010101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b00111101000110010100000110100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111110110000111000110001100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111101001010110100001000000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111101001110000110100000011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111110101100000000110001010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111101110001101111101110011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b10111110001100101010010100010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b00111110000001011000110111111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111100100100100010010100101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111100110100111011010001010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111101111001111100011110010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b10111101100001001100010111101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel6_Valid_Out)
	);
	Adder_64input add_k6(
		.Data1(Data_Out_Kernel6[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel6[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel6[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel6[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel6[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel6[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel6[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel6[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel6[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel6[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel6[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel6[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel6[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel6[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel6[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel6[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel6[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel6[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel6[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel6[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel6[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel6[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel6[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel6[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel6[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel6[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel6[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel6[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel6[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel6[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel6[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel6[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel6[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel6[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel6[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel6[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel6[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel6[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel6[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel6[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel6[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel6[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel6[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel6[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel6[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel6[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel6[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel6[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel6[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel6[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel6[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel6[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel6[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel6[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel6[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel6[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel6[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel6[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel6[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel6[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel6[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel6[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel6[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel6[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel6),
		.Data_Out(add_k6_Data_Out),
		.Valid_Out(add_kernel6_Valid_Out)
	);
	Batch_Norm bn_kernel6(
		.Data_A(32'b00111110010111100011001000001001),
		.Data_B(32'b10111110101100010101010000000001),
		.Data_In(add_k6_Data_Out),
		.Valid_In(add_kernel6_Valid_Out),
		.Data_Out(bn6_Data_Out),
		.Valid_Out(bn6_Valid_Out)
	);
	Relu_Core rl_kernel6(
		.Data_In(bn6_Data_Out),
		.Valid_In(bn6_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(rl6_Valid_Out)
	);
//////////KERNEL7//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111110110101111001010101010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110100010001100110011001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110110010010101010010010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110101101011001110111010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111101110001000100100101000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110100011100011100110101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111100101011110001100110110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111110011101001011000001100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110010110001111100011110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111100110011101111001101001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111100110100101111100111010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111110010111001101011101111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110010011100110011010010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111101110101100001101110011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110101001010000111010011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111110100011000100101010100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110010101010100010111000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111101100001011111000000110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111100110000011000001010101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110110100101010001010111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110101011110000110010101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111101101100010110011011111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111111000100100110101011110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111101100101000011101110100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111101110100001001001111111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110011111001000000110001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111101111011110011011010001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110110100000101010000000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111110100100010001110011000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111110010101111000000101111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111110001100011111111100000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110001110011001110010001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111111000001010101010110100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b00111110111000010010011101010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111111000001000000110111110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b10111110011011110000000101000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111110101010011001110110100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111101100001110100000011110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111101110100010101001111110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111100101101000001100011010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111110110100111000011010110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111110110010010100100010000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111110000001010100010010111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111101110000011011010101101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111110011110011111101010001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111110100011111101101000011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111110011110000110000100011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111110110101100001001101101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111110100011111101110100000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b00111110001011100010100100110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111110001011010110110110110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111110001011100101001011110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b00111101001000101001000100001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111110110011010101000000101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111101101000100011010000000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111101110011100100100101101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111110011100001101101110001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111011010111001101111110000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111010111000100011001101010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b00111101110010110010111110011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111110101100100100011100111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b10111101111010000100000111111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111100010111010000110111001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b10111101111101110011110010110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel7_Valid_Out)
	);
	Adder_64input add_k7(
		.Data1(Data_Out_Kernel7[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel7[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel7[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel7[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel7[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel7[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel7[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel7[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel7[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel7[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel7[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel7[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel7[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel7[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel7[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel7[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel7[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel7[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel7[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel7[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel7[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel7[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel7[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel7[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel7[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel7[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel7[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel7[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel7[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel7[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel7[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel7[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel7[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel7[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel7[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel7[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel7[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel7[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel7[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel7[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel7[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel7[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel7[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel7[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel7[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel7[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel7[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel7[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel7[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel7[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel7[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel7[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel7[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel7[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel7[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel7[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel7[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel7[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel7[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel7[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel7[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel7[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel7[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel7[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel7),
		.Data_Out(add_k7_Data_Out),
		.Valid_Out(add_kernel7_Valid_Out)
	);
	Batch_Norm bn_kernel7(
		.Data_A(32'b00111110010111010011111011110111),
		.Data_B(32'b10111110111100000011100001100001),
		.Data_In(add_k7_Data_Out),
		.Valid_In(add_kernel7_Valid_Out),
		.Data_Out(bn7_Data_Out),
		.Valid_Out(bn7_Valid_Out)
	);
	Relu_Core rl_kernel7(
		.Data_In(bn7_Data_Out),
		.Valid_In(bn7_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(rl7_Valid_Out)
	);
//////////KERNEL8//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111111000100000001000101100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110010000100101110010101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111100100110110111001011111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111101100011100001011101011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111110000110010101010010011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111101111000110111000101111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111110010100101010100000101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111100110100001101010010101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111101101000000001011101001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111101001110000110000010000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110000000110111101110001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111101101000110010101000101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110001000011111001010111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111101110110010010001101101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110010100010101010011000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111110010111011001011100110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110100001101110110000010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110000110001100000011000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110100100100110100100011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111101111100000001110000011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110011110000010011100111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111101101110111000000111001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110010010010000100000011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111101110100010111100100011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111101001010001111001010101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110110000011011100100101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110110100101001001010010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111101100110010010000000110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111101101101100100001111010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111110010101001000111111001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111110101101110011101010001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110010111001010011001100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b00111001011011000001000000001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b00111110100101010010111100001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111110101111001011000010110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111010010100001010010000001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111110100010101111001010010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111110010011000101000011011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111100001100111101001011101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111101111001101111101110000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111111001011011000110110110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111110010111111111110111011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111101111000100011101101001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111110010100011011100011010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111101110100101011101101100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111110101111011100011100101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111110110100001111001110011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111110000101111011111010000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b00111101001110001010101001010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b00111101000000110101111100101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111110000000001000001010000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111110000011100010110100111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111011110001111110010111001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111110110000010010011101000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111110010101011010001011001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111101100110010100111000100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111110101100011111011001001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111110011110000100101110000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b10111110001001011100000100010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b00111101000011010111001011110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111101001110001011001100011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111100100101111111110111000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111110110010010101010101001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b10111101000100111000101101100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel8_Valid_Out)
	);
	Adder_64input add_k8(
		.Data1(Data_Out_Kernel8[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel8[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel8[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel8[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel8[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel8[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel8[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel8[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel8[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel8[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel8[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel8[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel8[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel8[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel8[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel8[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel8[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel8[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel8[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel8[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel8[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel8[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel8[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel8[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel8[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel8[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel8[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel8[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel8[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel8[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel8[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel8[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel8[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel8[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel8[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel8[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel8[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel8[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel8[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel8[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel8[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel8[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel8[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel8[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel8[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel8[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel8[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel8[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel8[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel8[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel8[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel8[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel8[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel8[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel8[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel8[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel8[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel8[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel8[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel8[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel8[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel8[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel8[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel8[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel8),
		.Data_Out(add_k8_Data_Out),
		.Valid_Out(add_kernel8_Valid_Out)
	);
	Batch_Norm bn_kernel8(
		.Data_A(32'b00111110011010000100111111010001),
		.Data_B(32'b10111110101110111100100110100111),
		.Data_In(add_k8_Data_Out),
		.Valid_In(add_kernel8_Valid_Out),
		.Data_Out(bn8_Data_Out),
		.Valid_Out(bn8_Valid_Out)
	);
	Relu_Core rl_kernel8(
		.Data_In(bn8_Data_Out),
		.Valid_In(bn8_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(rl8_Valid_Out)
	);
//////////KERNEL9//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111111010111111011100100111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111110100010000011000000101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111101101000010011111100111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110010100010101001000110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111101000010110011100111110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110000110000011000101001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111110111100011100011000011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111101111011001010011011110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111110010010001111010010000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110011110000111001011100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111101001100110011011010001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111100000101111110000110000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111110111110011111001000010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111110110011001010010101010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110000110100011100101011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111101111011001000111001001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111101010000110001001100001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110010110101011110010101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110100100000111000010101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111101111100001100010010110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110111000000010100010110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111111010111100111101110001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110010001101100110110101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111110010101001000011111010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111110101100101101010111011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110011111101010111101101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111101111011001010011010000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111110100100010100011010010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111101111000011000110101101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111111001110000110101111010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111110001010011101000011101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110101011100011010001001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b00111111000111100001111011110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111110101110111010000110011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111110111100101011011010100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b10111110001011111110110110101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111101001010111010110111010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b00111110101111111111101111110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b00111111000110010100111000000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111110100111111010011011011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111110101011010010110001110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111110000011001001010110010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111110101111011011101101100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b00111110101010001011101001100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111110001110010011110010001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111110110111100111010111100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b10111110101010000000110101111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111110001011010010010010001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111110100100010010011010011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111110101100001111101011100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b10111101010100001101000000000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111110100111010101010100111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111100011111011010011101111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b00111100000010100110100001010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b10111111000000010000101001100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111101111011000000001001010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111111010010011010010110011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111101110010000101001111100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111110101110110001111010100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111110010000010001101100111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b10111100101001111000001110111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111110100100011101111000101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111101100000111011010111101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b10111110110000010100100000010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel9_Valid_Out)
	);
	Adder_64input add_k9(
		.Data1(Data_Out_Kernel9[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel9[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel9[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel9[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel9[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel9[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel9[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel9[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel9[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel9[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel9[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel9[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel9[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel9[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel9[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel9[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel9[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel9[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel9[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel9[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel9[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel9[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel9[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel9[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel9[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel9[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel9[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel9[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel9[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel9[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel9[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel9[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel9[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel9[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel9[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel9[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel9[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel9[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel9[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel9[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel9[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel9[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel9[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel9[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel9[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel9[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel9[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel9[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel9[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel9[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel9[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel9[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel9[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel9[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel9[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel9[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel9[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel9[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel9[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel9[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel9[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel9[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel9[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel9[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel9),
		.Data_Out(add_k9_Data_Out),
		.Valid_Out(add_kernel9_Valid_Out)
	);
	Batch_Norm bn_kernel9(
		.Data_A(32'b00111110010001111000011011110101),
		.Data_B(32'b10111110011011101101011001110010),
		.Data_In(add_k9_Data_Out),
		.Valid_In(add_kernel9_Valid_Out),
		.Data_Out(bn9_Data_Out),
		.Valid_Out(bn9_Valid_Out)
	);
	Relu_Core rl_kernel9(
		.Data_In(bn9_Data_Out),
		.Valid_In(bn9_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(rl9_Valid_Out)
	);
//////////KERNEL10//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110010101010011101001101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111110011011101111010101111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111101100011111000111001110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110101101101111111100110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111101010110100111110110111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111101100010100011001000110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111110110001001101001010011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111110000100101111101101111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111110011111101001111001011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111101010001110110100111010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111110000101110111110001001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110100001110001110011111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111011111000110010110100111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111101100100011111010000011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110110001000000110101011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111110001111100101100100100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111111001111101101001010000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111110000101000010110111101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111110011001010010101110010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111101110101010011111111111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110010111111000111000100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111101101001001000111001111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111110011111011111001001011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111110110001001110000100011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111101100110000111110000001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111110001001101111101111001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111110001101000101011010110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111101011000111110010101111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111100011001001000000100001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110111011010111100100101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111110001100011100100110100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111110101010001111000101010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b00111101101010111001101110111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111110010100110110011011011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111110010010100011011010110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111101101000001010101111010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b10111110101001001110101111000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b00111101100111001001011001001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111110111000000001011110101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b00111110100100000011100001000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b10111111010100100111010111010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111101101010000100011011111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b00111110010101100001010101111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b00111110000011011101111011111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b00111110101100111111110110010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b10111110001101001111111110111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b10111110110011101101100100000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b00111110100110110110001111100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b00111101010101000101101100111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111101000010000111100110110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111100101000001100011010000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b10111110100100101101011010111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111110000000111010011001001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b00111110001110011001011111001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111101110101111110000111100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111101110001000100101001001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b10111110011110100100100010100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b10111110101111011111100110101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111110000101110100011101110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111101001001100101010111111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111100100110100101000101100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111110001101000010100010110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b10111110101000110001100100101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111101110011001011111100011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel10_Valid_Out)
	);
	Adder_64input add_k10(
		.Data1(Data_Out_Kernel10[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel10[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel10[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel10[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel10[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel10[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel10[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel10[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel10[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel10[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel10[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel10[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel10[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel10[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel10[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel10[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel10[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel10[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel10[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel10[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel10[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel10[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel10[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel10[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel10[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel10[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel10[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel10[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel10[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel10[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel10[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel10[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel10[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel10[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel10[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel10[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel10[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel10[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel10[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel10[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel10[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel10[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel10[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel10[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel10[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel10[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel10[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel10[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel10[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel10[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel10[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel10[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel10[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel10[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel10[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel10[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel10[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel10[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel10[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel10[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel10[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel10[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel10[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel10[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel10),
		.Data_Out(add_k10_Data_Out),
		.Valid_Out(add_kernel10_Valid_Out)
	);
	Batch_Norm bn_kernel10(
		.Data_A(32'b00111110001010010101100011001110),
		.Data_B(32'b00111101000111001101111011000001),
		.Data_In(add_k10_Data_Out),
		.Valid_In(add_kernel10_Valid_Out),
		.Data_Out(bn10_Data_Out),
		.Valid_Out(bn10_Valid_Out)
	);
	Relu_Core rl_kernel10(
		.Data_In(bn10_Data_Out),
		.Valid_In(bn10_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(rl10_Valid_Out)
	);
//////////KERNEL11//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111111000010001100010101010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111110101010010010010100110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110010000100111001110011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111111000111000110101101100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111110101110000001011110001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110011101101010010110001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111110101011001110101100110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111101100000011101010111101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111110110101110101101010001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111110101111000110111100001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111101000001111110101010001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111111000010100011111010000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111101100011110100011001010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111110001100100110010001111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111011111010001100110101000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111110000101010010110001110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111110110010101111011100011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110100011011000111010110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110000001110101010111100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110111010001010111011000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111111011101010100011000011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111111001011000001110011100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111110010000010011110101001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111111000010011100001000100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111101011000110011111001011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111111000101100011010110001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111100110100111001100111110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111101100101111001100011101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111101100101101000110101000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111110010110010010110000011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111110111011111111100001000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111110001011001111000011000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b00111110111110010011110000110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111110111010111010111011100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111110100001111100100001011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b10111110100011111110001010101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b10111111001000011001111001110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b00111110101000110000101000101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111110001110011111011000111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b00111100110111101111000001101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b10111111000110010110000010010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b10111110100001010011101101101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111101100101110111011110110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b00111101100110101011100011001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b00111110100110011001011010010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b10111101101001110010001000101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b10111101100001001110111010101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111110010011010011010000111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111110011011111011100001110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111100110011010101100100011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b10111110000100011110100011011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111100110100111110010110011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111011101001100110110100001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b00111111010100001111111001000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111110001100011001101000000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111101011010000001111001010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111110010011000001110011010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111100000111111100000011000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111101100100010011101010000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b00111100000000101101001010001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b10111101111100100000000111100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111110111101101110111100011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b10111110101110001101000001011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111110000001001100010011101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel11_Valid_Out)
	);
	Adder_64input add_k11(
		.Data1(Data_Out_Kernel11[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel11[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel11[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel11[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel11[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel11[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel11[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel11[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel11[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel11[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel11[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel11[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel11[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel11[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel11[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel11[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel11[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel11[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel11[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel11[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel11[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel11[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel11[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel11[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel11[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel11[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel11[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel11[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel11[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel11[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel11[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel11[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel11[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel11[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel11[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel11[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel11[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel11[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel11[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel11[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel11[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel11[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel11[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel11[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel11[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel11[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel11[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel11[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel11[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel11[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel11[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel11[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel11[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel11[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel11[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel11[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel11[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel11[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel11[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel11[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel11[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel11[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel11[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel11[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel11),
		.Data_Out(add_k11_Data_Out),
		.Valid_Out(add_kernel11_Valid_Out)
	);
	Batch_Norm bn_kernel11(
		.Data_A(32'b00111110000110001001000101011101),
		.Data_B(32'b10111110000011101011111011111101),
		.Data_In(add_k11_Data_Out),
		.Valid_In(add_kernel11_Valid_Out),
		.Data_Out(bn11_Data_Out),
		.Valid_Out(bn11_Valid_Out)
	);
	Relu_Core rl_kernel11(
		.Data_In(bn11_Data_Out),
		.Valid_In(bn11_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(rl11_Valid_Out)
	);
//////////KERNEL12//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111111000101010001101011011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111100110010101101011100110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111111000100110010101011011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111111000101011000101101010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111110001111000001000000011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111110001010011000110101011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111110010110001000111001111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111110001000111110010110101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111100101111010101101010110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111110011111100111111010000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111111000110101010010111010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111110010010100001111010011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111101000111101100011111001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111110110111010001000010100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110100011101001011110110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111101001010010100101001011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111101001111101001110011100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110010011111000111111001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111111000110011100101011111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111101010010000011010000100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111101111000001110001000001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111101000110011011011001101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111111010001100111011011110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111110100100000010011001000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111111011111100000001111011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111111000001111011001110010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110001001011010110000000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111101110010000101011001011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111111000111100110110011010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110101101111111011110100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111101101100011110110000110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111101101100001010111111111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111011110110111000101000111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b00111101101100011010100101010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111110001101000000101101010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b10111110100101101011010101101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b10111111001100111101010001001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111110110011010101011011100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111111000100000010100110110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111110001101011010110101110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b10111110110110100110100001100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b10111110100111100100101011000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b00111110011111110101100001010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111111001001001111001110000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b00111110001100111010000010111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b10111101111111111001000110100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111110100001001010111001110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b00111100101001010001111011000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b00111110100010101101111010010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b00111110101111000010000010110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b10111110010001101001001000000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b10111110000010011111000000000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b00111101000110011001110111000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b00111110101000011011010011100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111101100000000101101000110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b00111101000010010110111101000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b10111111000100101000011110001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b10111110011110111110001001101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b10111110000001100100111101011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111100011011111001110101000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b10111110000110001000111001100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111101111101011111010100111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b10111110111000100010100100000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111110100110011011100010010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel12_Valid_Out)
	);
	Adder_64input add_k12(
		.Data1(Data_Out_Kernel12[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel12[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel12[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel12[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel12[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel12[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel12[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel12[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel12[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel12[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel12[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel12[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel12[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel12[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel12[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel12[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel12[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel12[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel12[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel12[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel12[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel12[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel12[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel12[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel12[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel12[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel12[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel12[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel12[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel12[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel12[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel12[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel12[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel12[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel12[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel12[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel12[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel12[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel12[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel12[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel12[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel12[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel12[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel12[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel12[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel12[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel12[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel12[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel12[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel12[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel12[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel12[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel12[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel12[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel12[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel12[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel12[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel12[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel12[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel12[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel12[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel12[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel12[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel12[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel12),
		.Data_Out(add_k12_Data_Out),
		.Valid_Out(add_kernel12_Valid_Out)
	);
	Batch_Norm bn_kernel12(
		.Data_A(32'b00111110001000001011101010001011),
		.Data_B(32'b00111111011110011011100010011100),
		.Data_In(add_k12_Data_Out),
		.Valid_In(add_kernel12_Valid_Out),
		.Data_Out(bn12_Data_Out),
		.Valid_Out(bn12_Valid_Out)
	);
	Relu_Core rl_kernel12(
		.Data_In(bn12_Data_Out),
		.Valid_In(bn12_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(rl12_Valid_Out)
	);
//////////KERNEL13//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110100001001010001001001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111110100111111000010011010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110100010110011000001111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110111100010110101011000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111101100011110110000000100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111101110110111111011010111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111101111000000001100000111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111100111110110000000001001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111110100111011011011100011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111100011001100000101111101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111100100000100000110010011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111101100101011111101111110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111100101001000010001111010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111101000010001100011001101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110100001100100000111001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111100111011101111111100111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111110111001111101010101110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110010010001101010000011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111101111100010001100011000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111101110100100110011101111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110110101001100000011011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111100001100101000000001000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111110101011110011001111000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111110101011110101010011011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111101000000110110010101111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111101110010011001100001111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111110101111101100001011110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111110100000000110011001100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111110100010100110101011010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110100110100000001100000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111101100010111110001010000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111110110101000101011101101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b00111110000000101011111001010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111101100110011110000010010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111101111111100110011111100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111110010000010001001011010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b10111110100101110110111010000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111110001011101101001101010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111110010001001101101110000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111101011001110100001001011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b10111111000100111110010110000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b10111100100101111011100111100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b00111110100011000101101101010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b00111101100011011001000110001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b00111110100000001110011111010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b10111110100110111111001111100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b10111101001001101110110011011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b00111110011100000100000010000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111101101011100111001011101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b00111101110111011001100000100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b10111101011100010000000010110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b10111110100100110000101101110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b00111101000101011011110110000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b00111110000101010011010011001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b10111100110110100001010001011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b00111101101110000111100010110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b10111110100101101100011000001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b10111110100010110000010010011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b10111100000010000111010110010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b00111100100001111100110001101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b10111110100001110100011111001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111110000100101011001010111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111101111000011111100000101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111101101110011011100110010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel13_Valid_Out)
	);
	Adder_64input add_k13(
		.Data1(Data_Out_Kernel13[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel13[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel13[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel13[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel13[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel13[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel13[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel13[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel13[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel13[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel13[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel13[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel13[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel13[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel13[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel13[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel13[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel13[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel13[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel13[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel13[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel13[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel13[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel13[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel13[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel13[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel13[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel13[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel13[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel13[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel13[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel13[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel13[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel13[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel13[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel13[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel13[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel13[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel13[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel13[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel13[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel13[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel13[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel13[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel13[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel13[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel13[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel13[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel13[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel13[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel13[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel13[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel13[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel13[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel13[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel13[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel13[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel13[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel13[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel13[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel13[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel13[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel13[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel13[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel13),
		.Data_Out(add_k13_Data_Out),
		.Valid_Out(add_kernel13_Valid_Out)
	);
	Batch_Norm bn_kernel13(
		.Data_A(32'b00111110010011100011101100010100),
		.Data_B(32'b00111111001100010010001011111000),
		.Data_In(add_k13_Data_Out),
		.Valid_In(add_kernel13_Valid_Out),
		.Data_Out(bn13_Data_Out),
		.Valid_Out(bn13_Valid_Out)
	);
	Relu_Core rl_kernel13(
		.Data_In(bn13_Data_Out),
		.Valid_In(bn13_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(rl13_Valid_Out)
	);
//////////KERNEL14//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111110101000101111010000001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110100001011001000000111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111101001010001101011101001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110110001010000111101101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111110011100011000001010101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110101000100101110100101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111110010010110110101010111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111101110111110010110110101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110010010101000010000100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110100000111100011000111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111101110110110011000001100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110010110001011010110110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110000010001101001010101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111101111010101101011110100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111101110111110000000100000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111110000100011100110011101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110001001101000000001100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111011011000101111100111110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111101110000011100001111000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111101100001101011011101010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111111000101111110100110011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111110011001011010100110111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111111000000111111111101110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111110101010110111100010011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111110110000000000100001001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111111010001011011000001000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111101110101001101001111011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111110010110000110010111100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111110111101101110110000101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111101000100111010101011111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111110001001000011010111000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111111010000101000110101100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111110110110011001011010011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111101111010000010001110110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111110010011100100100100010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111110100000110001001110101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111110110101011011001101101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b00111110000101011100101101011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b00111111000101011001101111010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111110011000000010010111010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111111010110101000011000100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111111001100100000101101101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111101110110000000110100111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b00111110101100010001010110111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111110100100001110110011111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111101011100001111011000101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b10111110001010101111100010011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111101100010100100101110001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111110100111110011001111100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111101110100011001011100001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111101101111000011101000111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111101011111111110011000010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111110010101011110010001000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111111001100101101101000110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b10111101110011000000010011001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b00111110001000101001000110110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b10111110001001110101000001001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111110010111000101001001110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111110010111010001110010101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111111001101011101011000011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111110110000010001101101110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111101101111110011010111110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111110111111111111100100000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b10111111000001010111001000010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel14_Valid_Out)
	);
	Adder_64input add_k14(
		.Data1(Data_Out_Kernel14[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel14[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel14[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel14[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel14[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel14[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel14[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel14[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel14[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel14[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel14[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel14[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel14[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel14[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel14[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel14[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel14[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel14[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel14[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel14[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel14[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel14[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel14[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel14[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel14[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel14[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel14[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel14[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel14[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel14[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel14[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel14[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel14[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel14[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel14[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel14[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel14[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel14[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel14[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel14[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel14[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel14[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel14[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel14[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel14[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel14[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel14[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel14[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel14[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel14[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel14[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel14[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel14[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel14[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel14[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel14[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel14[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel14[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel14[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel14[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel14[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel14[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel14[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel14[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel14),
		.Data_Out(add_k14_Data_Out),
		.Valid_Out(add_kernel14_Valid_Out)
	);
	Batch_Norm bn_kernel14(
		.Data_A(32'b00111110000101010000010010001011),
		.Data_B(32'b10111110101011010011001101100011),
		.Data_In(add_k14_Data_Out),
		.Valid_In(add_kernel14_Valid_Out),
		.Data_Out(bn14_Data_Out),
		.Valid_Out(bn14_Valid_Out)
	);
	Relu_Core rl_kernel14(
		.Data_In(bn14_Data_Out),
		.Valid_In(bn14_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(rl14_Valid_Out)
	);
//////////KERNEL15//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110010010010010110001111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111010110011001100011100001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111101010011110101100110100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111100101110010101000010100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111110010000110000100110000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110011101011100111011011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111101111111000110010010011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111101101111110110101110101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111101100000000010001101001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111101010000001110110011111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111101110011001110010000100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110000011001101101011100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111100100111111001101011111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111100110011111110100101000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110001111110010110100101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111111001011110001010011010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111110111111010100001101010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111101100100101010111001001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111110101101111110100011010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110000011110111111110010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110011111011110010110110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111101001100001010111010011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111100000110101000111011001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111110111101111100110101110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111110000010000111110011001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111110110110001111000101110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111111000010110000010110111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111101111000110000011101010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111100110000101000111011110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110110010101100110101110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111110011010100111011001100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111110011100111110111110110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b00111100000010001001101101010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111110100100000100010110010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111111010101101011010101000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111101111001100101110111100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111101001000010110101010111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b00111110001010010111101010111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111110101111110110001100101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b00111101000000110011010110011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b10111110110110111101011100011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111110010110101110000100110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b00111101101110101101100011111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b00111101100011110110010010001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b00111110110101100000000011010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b10111110101010001011010001000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b10111110000101001010000000101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b00111110101101111010100110111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111110000100000000001110011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b00111110010001110010000110000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111101111000101000011100001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b10111110100110001111000111100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111101100101001000001010100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b00111110100110001100010001010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111101000001001100101001011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b00111101111010101001110001101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b10111111000100100001011010001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b10111110001001111111110100011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111110010001111000011110010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b00111101011010001101100011001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111110100001100111000101011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111101111000011001011100000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b10111110000111000000101001111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111110000001001101101110100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel15_Valid_Out)
	);
	Adder_64input add_k15(
		.Data1(Data_Out_Kernel15[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel15[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel15[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel15[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel15[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel15[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel15[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel15[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel15[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel15[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel15[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel15[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel15[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel15[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel15[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel15[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel15[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel15[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel15[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel15[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel15[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel15[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel15[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel15[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel15[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel15[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel15[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel15[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel15[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel15[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel15[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel15[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel15[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel15[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel15[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel15[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel15[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel15[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel15[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel15[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel15[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel15[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel15[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel15[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel15[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel15[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel15[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel15[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel15[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel15[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel15[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel15[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel15[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel15[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel15[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel15[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel15[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel15[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel15[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel15[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel15[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel15[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel15[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel15[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel15),
		.Data_Out(add_k15_Data_Out),
		.Valid_Out(add_kernel15_Valid_Out)
	);
	Batch_Norm bn_kernel15(
		.Data_A(32'b00111110010011110011100010111110),
		.Data_B(32'b00111101101100000001100000101001),
		.Data_In(add_k15_Data_Out),
		.Valid_In(add_kernel15_Valid_Out),
		.Data_Out(bn15_Data_Out),
		.Valid_Out(bn15_Valid_Out)
	);
	Relu_Core rl_kernel15(
		.Data_In(bn15_Data_Out),
		.Valid_In(bn15_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(rl15_Valid_Out)
	);
//////////KERNEL16//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111111000001111000001010110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111110001010110011000000111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110000000001011000010010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110101001111010111011010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111101001111110011100001011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110010110111010111110000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111100001000010101101101011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111101101000110100001000101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110000101001011010111101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111101101100111110101111001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110011010010001010100110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111101110101011110010101100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111101101010001011110110111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111110100010101100101111000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110010001100101011111110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111110000101011100010100001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110000110101101101000001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110011001110110100010011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110011010111011001011001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111110001110001001011011110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110011110011101000000000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111110101101101000100010010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111111000000010111111111011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111111000110000101000111001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111110110000010000011100110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110101010011111001100000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110101001101110111101100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111110101111101000000100011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111110111000001100010110100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111111000000011010110110110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111101101010101000011011011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110101111110011011000100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111110100110111110111101011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111110001001000011000111010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111110000111111110111100000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111101110100101000100100101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111110001110001010001000000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b00111110001111010111000100010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b00111111001011101100110101101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111110110010100011011100101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111111011101000110010100101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111110100111101111010101001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111110011011100100111000101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b00111111000010000011110001101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111110110001101011000111111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111110001110011101010100110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b10111110010011110000001110000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111110010001101111111000000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111110100010100011011111001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111101100100111100001101000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111110101010010110010100111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111110011111011000011001001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111101010010011011111100111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111111001011101001100101111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111110000100000001101101100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b00111101100111111111111110010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111110101011110100111001100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111110101010010101110010011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111101100100010010001001010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111110111110100111110011110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111110101101111111110110100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111101111111100001000000100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111111000110111011000001110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b10111110110101110011111000101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel16_Valid_Out)
	);
	Adder_64input add_k16(
		.Data1(Data_Out_Kernel16[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel16[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel16[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel16[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel16[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel16[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel16[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel16[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel16[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel16[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel16[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel16[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel16[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel16[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel16[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel16[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel16[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel16[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel16[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel16[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel16[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel16[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel16[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel16[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel16[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel16[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel16[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel16[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel16[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel16[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel16[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel16[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel16[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel16[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel16[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel16[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel16[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel16[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel16[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel16[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel16[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel16[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel16[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel16[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel16[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel16[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel16[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel16[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel16[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel16[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel16[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel16[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel16[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel16[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel16[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel16[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel16[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel16[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel16[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel16[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel16[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel16[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel16[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel16[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel16),
		.Data_Out(add_k16_Data_Out),
		.Valid_Out(add_kernel16_Valid_Out)
	);
	Batch_Norm bn_kernel16(
		.Data_A(32'b00111110000011001001010101010110),
		.Data_B(32'b10111110101111101110110100010010),
		.Data_In(add_k16_Data_Out),
		.Valid_In(add_kernel16_Valid_Out),
		.Data_Out(bn16_Data_Out),
		.Valid_Out(bn16_Valid_Out)
	);
	Relu_Core rl_kernel16(
		.Data_In(bn16_Data_Out),
		.Valid_In(bn16_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(rl16_Valid_Out)
	);
//////////KERNEL17//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110011101110010001101011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111110010110000010010110100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110000011001011100011110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110100010011110100101100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111101010011010110101110101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110000101000110011011111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111110011111000100101011001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111011110101011110011010110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111110111110111001011110100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110001110001100001011001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111101111000010111100100100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111101001000010000010110001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111010101101000110011000100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111110101100100101001101101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110100101110100000110110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111110010110111111111110001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111110011001001101100011100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111110001010010010001010101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111101100010110110110010001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111101100001100110011110110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110110000111001011100010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111110000010110011101001101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111110010111110110011001000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111110100111011000101101111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111101100100111011010001110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111110001010001000101101111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111110111001011010101000101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111111000010101110001001111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111101100010011100101110010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110110110110010111010111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111110011001011100001010001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111101100000001000011001011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b00111110011000100000000101111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111110100101101010000000001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111111001100001001001100010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111110010010101111101101101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b10111101101000101100101111000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b00111110001101100001111000101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111110111001001100111100110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b00111101001110111101000100110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b10111110110101000111111101010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111110001010101100100011011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b00111110001001100011001100100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111101010011100100110011101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b00111110111011100000100100011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b10111110011000111101111100110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b10111110001000100000010111011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b00111110110101100110111000100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b00111101100001010011011111000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b00111110011110110010001100101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111110010000000010011110011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b10111110100111000011001100010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111110010010010011100011100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b00111110010001111010000000001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b10111110000100101000001101010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b00111110001000000111111100101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b10111110111001001100100110011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b10111111000111111100011100100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111110101011111000111110101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111110000111100001111101001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111101111101101000110011111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111110010001101000000111111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b10111101101101101110010010011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111101001010001001011111100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel17_Valid_Out)
	);
	Adder_64input add_k17(
		.Data1(Data_Out_Kernel17[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel17[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel17[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel17[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel17[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel17[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel17[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel17[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel17[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel17[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel17[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel17[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel17[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel17[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel17[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel17[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel17[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel17[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel17[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel17[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel17[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel17[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel17[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel17[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel17[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel17[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel17[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel17[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel17[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel17[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel17[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel17[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel17[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel17[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel17[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel17[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel17[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel17[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel17[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel17[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel17[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel17[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel17[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel17[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel17[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel17[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel17[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel17[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel17[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel17[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel17[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel17[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel17[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel17[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel17[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel17[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel17[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel17[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel17[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel17[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel17[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel17[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel17[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel17[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel17),
		.Data_Out(add_k17_Data_Out),
		.Valid_Out(add_kernel17_Valid_Out)
	);
	Batch_Norm bn_kernel17(
		.Data_A(32'b00111110001111010000010011011001),
		.Data_B(32'b10111110100100010011010010110001),
		.Data_In(add_k17_Data_Out),
		.Valid_In(add_kernel17_Valid_Out),
		.Data_Out(bn17_Data_Out),
		.Valid_Out(bn17_Valid_Out)
	);
	Relu_Core rl_kernel17(
		.Data_In(bn17_Data_Out),
		.Valid_In(bn17_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(rl17_Valid_Out)
	);
//////////KERNEL18//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111111000110011011010000010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111110001001001000101001100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110010110010110101010110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110010101100010111111100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111101100011101100100110111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111101011101010001110100111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111110000100000011001110110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111100100111010011100000110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110100110000000000111101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111100110011100001001001101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111101100011100001100101000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111110100001010111111000100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110011001010011101001010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111101111001010011000010001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110010001101111101011101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111110001001101010101010110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111111000001111010000011100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111101110010001110010011110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111101111100111001100010000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110100101011011000110110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110001101001010011011000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111101100100001100101000110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110101101011001100011100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111101101111111000101000100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111110111001110110101000001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110010000101101100110110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110001011101110011100000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111101101111101001001010111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111110000001001101101010100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111101001000110101010110001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111101101110011110010001111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111101010100010001111111101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111110001110101111101101000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b00111110011111110000010111101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111111000000101111001000000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b10111100100101101001101000110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111110110110010100000101011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111110000001110100001111101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b00111101111100110101111111110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111110010011100100111010001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111110110000111010100001010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111110000101000001010111011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111101100001010101110111000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111101010111010101100011000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111101101011110001010000010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111110011001110110101001100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111110110001010110000111010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111110110010011010110000101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111101001111110111101110010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111101001100101110110001110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111101000110100001011011110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111110000110101010010111010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b00111101101011110110000011100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111110111010011101010101000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b10111101010001011111101110110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111101110110111100110110001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111110101000110011001110100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111100110000010010110010001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b10111110001100110000000010001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b00111110000011110110110001101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111101001111000001100000110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b10111101101010111001011000111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b10111101110101100001010010101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b10111101100111100101100111011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel18_Valid_Out)
	);
	Adder_64input add_k18(
		.Data1(Data_Out_Kernel18[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel18[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel18[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel18[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel18[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel18[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel18[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel18[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel18[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel18[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel18[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel18[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel18[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel18[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel18[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel18[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel18[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel18[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel18[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel18[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel18[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel18[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel18[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel18[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel18[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel18[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel18[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel18[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel18[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel18[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel18[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel18[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel18[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel18[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel18[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel18[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel18[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel18[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel18[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel18[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel18[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel18[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel18[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel18[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel18[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel18[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel18[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel18[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel18[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel18[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel18[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel18[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel18[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel18[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel18[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel18[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel18[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel18[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel18[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel18[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel18[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel18[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel18[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel18[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel18),
		.Data_Out(add_k18_Data_Out),
		.Valid_Out(add_kernel18_Valid_Out)
	);
	Batch_Norm bn_kernel18(
		.Data_A(32'b00111110010111100110100100111000),
		.Data_B(32'b10111110100111101101010111001110),
		.Data_In(add_k18_Data_Out),
		.Valid_In(add_kernel18_Valid_Out),
		.Data_Out(bn18_Data_Out),
		.Valid_Out(bn18_Valid_Out)
	);
	Relu_Core rl_kernel18(
		.Data_In(bn18_Data_Out),
		.Valid_In(bn18_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(rl18_Valid_Out)
	);
//////////KERNEL19//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111111000100010101111000110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111101101010011001100111110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110011011101011100111111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111111000001100000101101100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111110001101101111111101110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110010111000001100110001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111101100101001111001100000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111110001001110100011011011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110100101011110001110011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110000011111001100000001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111101111000010001000111101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111110100000110110111010000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110010100101001011000001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111101010110011010011001110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110101100001001111100010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111101101101011011100011001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110110010110111100010000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111010011000010000100111011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110100000101100111001111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110110101111010001100001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110010011011110000011010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111101101111000010111110001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110110101100101011101001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111101101001001101101110000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111110110011111010111110111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110000010111110110011001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111101001000111010000100000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111010111110111100011111100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111110000110011010110000001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111110100111010110110101000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111110001100000101111101111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111101100101100001000001011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111110000001111011111000101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b00111101101001111110001010011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111110110001000010001100100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b10111010100010100110111100100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111110101000000011011111001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b00111100011111001101101111001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b00111101101101000111001101101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111101111010000000011101011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111111000010111011010001111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111110011110000001011111111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111110010000011011110110011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111110010110100000101010011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111101101000111101100101000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111101100001010111101010000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111110011101010000110011100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111110110001010001011001000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111110000101011100110111011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111100101101111001010100101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111110100001011001111111001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111101111111010111101110110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111100011100111001110000001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111110101101100111000101111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111101000001110111010000000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b00111101100100111011111010000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111110001110100100100101111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111101000011010111011110100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111101000110111001111010001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111101101001110000011101000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111110001100101001011110101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111100001011000110101000100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111110000000011000000001011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b10111110000101010111001010000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel19_Valid_Out)
	);
	Adder_64input add_k19(
		.Data1(Data_Out_Kernel19[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel19[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel19[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel19[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel19[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel19[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel19[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel19[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel19[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel19[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel19[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel19[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel19[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel19[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel19[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel19[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel19[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel19[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel19[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel19[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel19[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel19[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel19[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel19[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel19[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel19[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel19[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel19[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel19[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel19[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel19[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel19[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel19[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel19[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel19[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel19[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel19[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel19[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel19[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel19[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel19[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel19[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel19[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel19[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel19[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel19[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel19[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel19[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel19[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel19[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel19[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel19[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel19[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel19[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel19[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel19[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel19[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel19[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel19[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel19[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel19[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel19[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel19[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel19[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel19),
		.Data_Out(add_k19_Data_Out),
		.Valid_Out(add_kernel19_Valid_Out)
	);
	Batch_Norm bn_kernel19(
		.Data_A(32'b00111110011001010001000111001110),
		.Data_B(32'b10111110100000101110011010111011),
		.Data_In(add_k19_Data_Out),
		.Valid_In(add_kernel19_Valid_Out),
		.Data_Out(bn19_Data_Out),
		.Valid_Out(bn19_Valid_Out)
	);
	Relu_Core rl_kernel19(
		.Data_In(bn19_Data_Out),
		.Valid_In(bn19_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(rl19_Valid_Out)
	);
//////////KERNEL20//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110100000001101001101101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111101111011110011110001101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110101100110111100000000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111101001110001101010011100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111110001110111000110001000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111110010011100010110100111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111111001111001000010000100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111110101000100001010011100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111100111000001111011010110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110111101101001111001000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111101100011011000010011100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110110100111001001101000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110100010001100000000101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111110010010000001110111010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110100001100101001101101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111111000111110111100001100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111110110101011000100101101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110000101100101100111100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110101011100011000011100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110000111010111000000110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110100101011101100001110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111110100000010001101100100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111110011011100110011111111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111110100001100011011100101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111111001010001010101000010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110010111101011000100101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111110110011000100100010100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111101100000100101111110000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111110101000001100111010111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111111001100010111111101000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111110010011110010001101011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111110100010101010110011011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b00111110100011111110111011101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111110110000000001000110111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111111001000100010001100111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111101111111010001000101100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b10111111000101110010111100010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111111000000011100001110101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111110100110001111101100010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b00111110101101000010000010110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111110000110010000110100010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111100101011000110100110111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111101001010101011111111000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111110101010010110001101000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b00111110101001001000110000111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b10111110010011100111011011001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111101101101011111101110001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b00111110010101110001011110000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b00111110111011010101100010100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111101001100100000101010101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b10111110001000001001100111100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b10111110100110110100001011101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111111001101101111001111100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b00111101100110010011111101100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111110100110000000000101110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b00111110001100101111000000101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b10111111001111001000010101011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111101001111110011111111110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111101100111110001110000110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b00111110001001100011111011100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111101110101010100011110101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111110011100011110101100010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111110001101001001100111100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b10111110110011011010010010011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel20_Valid_Out)
	);
	Adder_64input add_k20(
		.Data1(Data_Out_Kernel20[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel20[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel20[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel20[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel20[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel20[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel20[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel20[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel20[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel20[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel20[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel20[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel20[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel20[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel20[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel20[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel20[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel20[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel20[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel20[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel20[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel20[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel20[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel20[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel20[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel20[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel20[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel20[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel20[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel20[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel20[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel20[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel20[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel20[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel20[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel20[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel20[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel20[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel20[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel20[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel20[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel20[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel20[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel20[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel20[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel20[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel20[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel20[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel20[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel20[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel20[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel20[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel20[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel20[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel20[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel20[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel20[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel20[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel20[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel20[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel20[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel20[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel20[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel20[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel20),
		.Data_Out(add_k20_Data_Out),
		.Valid_Out(add_kernel20_Valid_Out)
	);
	Batch_Norm bn_kernel20(
		.Data_A(32'b00111110000100110001010100111011),
		.Data_B(32'b00111101110110111001001110001110),
		.Data_In(add_k20_Data_Out),
		.Valid_In(add_kernel20_Valid_Out),
		.Data_Out(bn20_Data_Out),
		.Valid_Out(bn20_Valid_Out)
	);
	Relu_Core rl_kernel20(
		.Data_In(bn20_Data_Out),
		.Valid_In(bn20_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(rl20_Valid_Out)
	);
//////////KERNEL21//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111111001010010101101011011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111101100010101110100101000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110010011101111100010001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110110100100110000111001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111100100100100110100011010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110001111101001001111001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111101000000110100011101010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111100110101100101001011111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110001010110001011101010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110000101000001100110010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110001100001111100100011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111101100000111110001100101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110000001100100111100111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111101111101111110000110000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111101101100010001110001001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111110010011011100111111110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111101110000010001111001001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110100110010011011010010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110100100110001011001101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111101100001100010000101100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110100001110100110100110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111110011111011001010010011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111111000100000001101000000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111110100001000100100000101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111100000101111011001100110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110001110111111101111111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110110000001011111110101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111101111011011001000010001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111101011011010010000101101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111111010011011011100000110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111101111101001011110101101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110011110101010010100000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111110010100111101011010110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111101001000011110000010101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111110110000001110100111011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b10111101101101111101101010100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111110001100110010011101011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111110010000001011101110110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b00111110100110100000101000011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111110100110111001001011011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111111001011011101011010001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111110010111000001100010001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111110011101001110010100001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111101000001011110110000101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111110111011010101111101001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111110100100011000000110110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111100010001011010101101111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111101110100000110110011100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111110001101011110110001101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111110010001111010110101111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111111000011111010111011000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111110100000000001010111011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111101010100001100010010110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111110100010000001011100100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111111000111100000001010011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111101001011110100100110011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111101100110111000110000111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111110110011101001110010110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111110000101111000010000111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111110010110110010011111110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111110100000010100000101110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111110100110101110101101111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111111000100111011011000000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b10111110010101001010001000110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel21_Valid_Out)
	);
	Adder_64input add_k21(
		.Data1(Data_Out_Kernel21[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel21[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel21[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel21[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel21[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel21[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel21[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel21[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel21[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel21[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel21[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel21[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel21[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel21[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel21[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel21[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel21[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel21[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel21[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel21[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel21[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel21[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel21[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel21[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel21[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel21[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel21[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel21[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel21[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel21[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel21[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel21[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel21[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel21[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel21[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel21[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel21[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel21[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel21[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel21[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel21[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel21[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel21[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel21[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel21[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel21[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel21[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel21[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel21[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel21[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel21[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel21[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel21[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel21[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel21[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel21[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel21[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel21[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel21[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel21[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel21[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel21[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel21[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel21[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel21),
		.Data_Out(add_k21_Data_Out),
		.Valid_Out(add_kernel21_Valid_Out)
	);
	Batch_Norm bn_kernel21(
		.Data_A(32'b00111110001111100100011110101000),
		.Data_B(32'b10111110110100100110010111100010),
		.Data_In(add_k21_Data_Out),
		.Valid_In(add_kernel21_Valid_Out),
		.Data_Out(bn21_Data_Out),
		.Valid_Out(bn21_Valid_Out)
	);
	Relu_Core rl_kernel21(
		.Data_In(bn21_Data_Out),
		.Valid_In(bn21_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(rl21_Valid_Out)
	);
//////////KERNEL22//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111101101000010001010110011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111101111000110000110000110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110001101010011110101110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111111000101010001011000100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111101011000010011101101100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111101010110111000100110001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111101111101010111111001111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111011111000000110010111110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111101100110010000101001101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111101101101010001000100110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111100011010111011000001001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110100000110100001001101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111100001000011011010110111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111100001111001100001010011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110101000101010100011101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111110010010001001100011011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111111011101110010010100101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111010110111110110100101010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111110010000111110111111010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111110011011110110100000000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110001000010001110001010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111110010011001101010010011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111101010111110100001110000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111110111110111101011000001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111101110110000110001101100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111110001101100100011100100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111101110000010101011100110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111100011010001101101000101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111110011010110100101111000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110001010111100110011010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111101111101100100110100011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111110101011000101110111011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b00111110000011101010110101110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111101110011100011111010010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111110110000010100000000001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111110011010011000111010110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b10111110010011001001010100101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111101100001011101111110011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111111000111001111000011111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b00111110100110000110010111101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b10111110101111111011010010100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111110001100101100100000111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b00111011000101101001111011001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b00111101100111100011110011011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b00111110100110011111011010010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b10111110010000101010100101101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b10111100110010100010110011001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b00111110100110001010101011001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b00111101110111001101000111111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111011111111101110110000101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b10111110000101001000100100001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b10111110111011000000010111110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111110100001001111100111100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b00111110100011111011101101000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111110011101010100011101001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b00111011101101110111001001010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b10111110111101111100110111000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b10111100101001011001001011011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b10111101011000001001001011111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b00111011111111000010011110111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b10111101111001101011100011110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111110000110101101101100000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111110001101010110011011011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111110010111001100010001001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel22_Valid_Out)
	);
	Adder_64input add_k22(
		.Data1(Data_Out_Kernel22[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel22[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel22[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel22[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel22[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel22[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel22[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel22[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel22[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel22[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel22[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel22[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel22[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel22[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel22[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel22[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel22[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel22[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel22[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel22[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel22[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel22[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel22[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel22[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel22[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel22[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel22[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel22[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel22[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel22[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel22[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel22[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel22[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel22[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel22[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel22[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel22[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel22[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel22[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel22[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel22[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel22[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel22[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel22[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel22[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel22[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel22[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel22[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel22[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel22[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel22[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel22[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel22[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel22[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel22[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel22[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel22[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel22[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel22[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel22[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel22[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel22[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel22[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel22[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel22),
		.Data_Out(add_k22_Data_Out),
		.Valid_Out(add_kernel22_Valid_Out)
	);
	Batch_Norm bn_kernel22(
		.Data_A(32'b00111110001111100111111001010101),
		.Data_B(32'b00111111000100011011011011010001),
		.Data_In(add_k22_Data_Out),
		.Valid_In(add_kernel22_Valid_Out),
		.Data_Out(bn22_Data_Out),
		.Valid_Out(bn22_Valid_Out)
	);
	Relu_Core rl_kernel22(
		.Data_In(bn22_Data_Out),
		.Valid_In(bn22_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(rl22_Valid_Out)
	);
//////////KERNEL23//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111110110100001100101110110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110001110110011101011100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110100101010110100110000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110011110000111111101111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111101110101101100010101010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111101101111001011001110101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111101111110011001111101110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111101110001110101111101001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111101101011101100000011111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111101101101101010110000100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110001001010101101110100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111101110000110111100101011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111011101001110111000001110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111110000000111110001000110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110000111001100111100001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111110000100111011001011100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111101101000001110111010100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111101101010011000001111010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111100110100101011111101000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111101101100011011001101110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110110000010001110000100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111100111001011001010001110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110100000110110111001101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111101101101110100100011000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111101101011001010111001100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110101010110100011011101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110111110100010011100111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111101110100101110110111111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111110100110101011101110011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111101110010100011100101100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111110101110011100001110001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110100011011010111100001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111110010010001100110011001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b00111110011001000101000100000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111110111111110101000010001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b10111110000111000110111011111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111110101100000110100111001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111110010001011101010001100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111100111111111111110000000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111101111111000010110101100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111111000101011000011111100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111110011010001100001001011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b00111101100100001110011010010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111101101101000100001000110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111101100000100101000110111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111110100010110000010110001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111101101111001100100100111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111110010010001000101000010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111101000110101000100001100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b00111101011011110110111011001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111110000100101100000000011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111100111101111000010111000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b00111110100000001111000011010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111110110011110011010000000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111110001000011110011111010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111110010011101110001011101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111110110000011010000110001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111110000101010010011101110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b10111101101010110100110111011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b00111110001100011000100101001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111101010000000100101110111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111101101100101110001111000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111110000111101001111111110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b10111100111110101001011100100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel23_Valid_Out)
	);
	Adder_64input add_k23(
		.Data1(Data_Out_Kernel23[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel23[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel23[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel23[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel23[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel23[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel23[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel23[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel23[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel23[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel23[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel23[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel23[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel23[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel23[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel23[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel23[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel23[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel23[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel23[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel23[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel23[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel23[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel23[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel23[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel23[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel23[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel23[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel23[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel23[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel23[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel23[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel23[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel23[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel23[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel23[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel23[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel23[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel23[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel23[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel23[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel23[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel23[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel23[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel23[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel23[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel23[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel23[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel23[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel23[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel23[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel23[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel23[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel23[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel23[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel23[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel23[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel23[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel23[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel23[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel23[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel23[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel23[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel23[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel23),
		.Data_Out(add_k23_Data_Out),
		.Valid_Out(add_kernel23_Valid_Out)
	);
	Batch_Norm bn_kernel23(
		.Data_A(32'b00111110011001101100000111001000),
		.Data_B(32'b10111111001011011011100111110000),
		.Data_In(add_k23_Data_Out),
		.Valid_In(add_kernel23_Valid_Out),
		.Data_Out(bn23_Data_Out),
		.Valid_Out(bn23_Valid_Out)
	);
	Relu_Core rl_kernel23(
		.Data_In(bn23_Data_Out),
		.Valid_In(bn23_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(rl23_Valid_Out)
	);
//////////KERNEL24//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111111000101100010110111001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111101010011110000010101010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110101011010111000100111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110111000111010101110010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111101111111000010101111000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111101110111110011100110100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111101101010110110011000101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111101111010110000001100000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110010011000001101000010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111100110001010000001101001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111110000000000100011100010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111110100010011110100100000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110100110100101011101000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111101111111011010000110100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110101010010010011001101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111110000100001000010000100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111111000110100110111111000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111110001001011001110001011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111101001111000100100110111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110101100000111101011110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111101100111010100010001110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111110001001010011000111010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110100110011110111100100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111101001000010111100101000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111110110101101010001001110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110000001101001000111001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111101101000101100100110110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111101100001100110111010111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111110010001101011110010110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110011010111000110101101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111110011011100001011100001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111101011011100001110100110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111110100111111001100111000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b00111101000011110010010010000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111110101100110100011010101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b10111101010100100010000110111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111110111000110000011001100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b00111101100000110101110010010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b00111110010011111011010110010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111101111000001110010000011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111110001111010110010000011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111110010110011000011010111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111101010001010000100011100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b00111110001000000101001101000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111110010011011101001001010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111011100110011001110011011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111110100010010100100110101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111110100011000101100110001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111110000100100101111000110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111101111001011100101011100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111110000100011110011001001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111110000000100000100010111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b00111100110100010010100000101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111110111001110100001010011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111100110100101111011111101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b00111110001011111001001111011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111110101000011000000011101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111101000100100011100100010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111110000100111110110100010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b00111110000010101010101000010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111110100011011100101010010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b10111101100011101101011001010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b10111110011001011011000001111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111110010011101101111010011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel24_Valid_Out)
	);
	Adder_64input add_k24(
		.Data1(Data_Out_Kernel24[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel24[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel24[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel24[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel24[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel24[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel24[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel24[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel24[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel24[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel24[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel24[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel24[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel24[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel24[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel24[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel24[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel24[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel24[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel24[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel24[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel24[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel24[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel24[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel24[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel24[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel24[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel24[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel24[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel24[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel24[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel24[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel24[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel24[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel24[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel24[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel24[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel24[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel24[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel24[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel24[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel24[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel24[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel24[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel24[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel24[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel24[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel24[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel24[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel24[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel24[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel24[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel24[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel24[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel24[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel24[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel24[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel24[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel24[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel24[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel24[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel24[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel24[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel24[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel24),
		.Data_Out(add_k24_Data_Out),
		.Valid_Out(add_kernel24_Valid_Out)
	);
	Batch_Norm bn_kernel24(
		.Data_A(32'b00111110011100011101011000111101),
		.Data_B(32'b10111111011000010001101001101010),
		.Data_In(add_k24_Data_Out),
		.Valid_In(add_kernel24_Valid_Out),
		.Data_Out(bn24_Data_Out),
		.Valid_Out(bn24_Valid_Out)
	);
	Relu_Core rl_kernel24(
		.Data_In(bn24_Data_Out),
		.Valid_In(bn24_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(rl24_Valid_Out)
	);
//////////KERNEL25//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111110001011111101101111110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110100101000111010101000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110001011011010101011001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110100011110011010111101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111110100010111100001110010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110000000110101000001100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111110101010110101000010010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111101000001000000101000100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111111010111001001101111011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111011100010000000101001101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110101001100101101001111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111110000111011101000111010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110011001000011111101011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111110000011001110001110011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111101100111101101000011100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111110000010100110000001011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110101011001101110011110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111101100111001111000001101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111110010000011100010100111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110010111010010001011111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110111100000001001011001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111110011001010011010001111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111101101111100000001110010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111111001101001101111011000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111110001111000110001111110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111101010101000011110110100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111111001101010100111000110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110100010100011100100010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111110010101111110110101000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110010001110111100110011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111110110110001001001001000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111100100001010110101100001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111111000110101100000110001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b00111110111100110111001110011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111110110000111001000001100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b10111100111000010101001000000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111111000011100110010001011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111110101111101111101001100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b00111101110011111111100110100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b00111101110010100001101101011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111111001100001010010101000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b10111100101010011100100010011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111110001001001101110111001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111101010000010110000110001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111110110101111100001001110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111111000110111111000010011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111110000111001001100010001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111110111110011110100110011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111110010100110111000010100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111101101000110111101011110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111011001010110010100100001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111110101101101100101111100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111110011010101111010110100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111111000110001001110000101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111010110011011010100010100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111111000111010001010111011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111101111111011110110010101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111110000111110010101101110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b10111110001001001010101101101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b00111110101001010101001000000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b10111101001010110100010101011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111110010001111100101111011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b10111110001001111000100100101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111110000011011010100011000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel25_Valid_Out)
	);
	Adder_64input add_k25(
		.Data1(Data_Out_Kernel25[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel25[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel25[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel25[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel25[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel25[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel25[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel25[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel25[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel25[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel25[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel25[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel25[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel25[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel25[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel25[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel25[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel25[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel25[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel25[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel25[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel25[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel25[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel25[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel25[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel25[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel25[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel25[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel25[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel25[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel25[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel25[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel25[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel25[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel25[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel25[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel25[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel25[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel25[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel25[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel25[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel25[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel25[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel25[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel25[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel25[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel25[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel25[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel25[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel25[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel25[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel25[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel25[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel25[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel25[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel25[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel25[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel25[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel25[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel25[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel25[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel25[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel25[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel25[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel25),
		.Data_Out(add_k25_Data_Out),
		.Valid_Out(add_kernel25_Valid_Out)
	);
	Batch_Norm bn_kernel25(
		.Data_A(32'b00111110000011101010000101010111),
		.Data_B(32'b00111110010000111101111000111100),
		.Data_In(add_k25_Data_Out),
		.Valid_In(add_kernel25_Valid_Out),
		.Data_Out(bn25_Data_Out),
		.Valid_Out(bn25_Valid_Out)
	);
	Relu_Core rl_kernel25(
		.Data_In(bn25_Data_Out),
		.Valid_In(bn25_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(rl25_Valid_Out)
	);
//////////KERNEL26//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110110011100000110010110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111110101111100111011101001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110000010011001101000100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110101101111001000100011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111101110101100010010101101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111010101010100110101010011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111110001111100101010101001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111110100010101001010110100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111110101111100000100101111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110010011101011111000000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111101011000110100000110110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110010001010110010111000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111101000011101110111101110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111101011001110011101010000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110111101010000001000011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111101110011011111101101000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111110101110010011100100101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111110000010110111101000110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111110000000010101100111010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111110001101000101110110110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110100100101011010010110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111110000111010000100111100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111110110110100101101111011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111110000111011000111110001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111101111001101111110110111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111110000111011010010100110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111110100100101000101011111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111110110100100000111101000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111100001000100111011111011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111111000100100100001100101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111010100000010011000100011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111110100001110110101001110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b00111100111011010010101000011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111110101110000000001011001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111110111011101100100110110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111110000011101100101101100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b10111101110000010001110100011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111110000111111110011100100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111110100101101010100000000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111101101001101100000101100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b10111111000011001100110010001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b10111100011011010110100100101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b00111110000101000101100101100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b00111101110111011110010001011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b00111110000001010100011111000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b10111110100001000111101010000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b10111110000111110000011101111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b00111110110111101111001001101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b00111101100111011100000010110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b00111101010100000100010110010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b10111100101100110101100100100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b10111110100001110110110101000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111101101101011110001001011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b00111100101100110111110001010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111110001001111000100011100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111100011100011100000110110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b10111101101110111100110001101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b10111110100101111001001000110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111110011110011010101111110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b00111110001001000110100000110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b10111100000011001000001100011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111101000001110011010001110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111100100010011111100001100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111110110001111001001000000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel26_Valid_Out)
	);
	Adder_64input add_k26(
		.Data1(Data_Out_Kernel26[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel26[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel26[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel26[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel26[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel26[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel26[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel26[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel26[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel26[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel26[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel26[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel26[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel26[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel26[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel26[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel26[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel26[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel26[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel26[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel26[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel26[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel26[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel26[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel26[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel26[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel26[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel26[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel26[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel26[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel26[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel26[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel26[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel26[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel26[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel26[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel26[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel26[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel26[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel26[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel26[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel26[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel26[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel26[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel26[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel26[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel26[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel26[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel26[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel26[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel26[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel26[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel26[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel26[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel26[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel26[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel26[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel26[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel26[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel26[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel26[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel26[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel26[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel26[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel26),
		.Data_Out(add_k26_Data_Out),
		.Valid_Out(add_kernel26_Valid_Out)
	);
	Batch_Norm bn_kernel26(
		.Data_A(32'b00111110010101111010001011100011),
		.Data_B(32'b00111101011011101011000011100000),
		.Data_In(add_k26_Data_Out),
		.Valid_In(add_kernel26_Valid_Out),
		.Data_Out(bn26_Data_Out),
		.Valid_Out(bn26_Valid_Out)
	);
	Relu_Core rl_kernel26(
		.Data_In(bn26_Data_Out),
		.Valid_In(bn26_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(rl26_Valid_Out)
	);
//////////KERNEL27//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111110101100001110001001110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110000000100111000110111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110000111101011010110001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110000110000101101000001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111100011001111000001000011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110000001101011011100100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111110011101100110001011000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111101101001000101111111010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111111000000101011001101100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111110010101010001001011001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110001001000001010100010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111101100101100010010011111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111101111001101010110011010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111110010010111101011000100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111101100101011011101001011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111110000111100000110111100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110100110001000100011010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111101101101000101000010100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111110010001101100000000011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110110011110100001000011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110101011101100010010000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111110000100101100111110011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110011100001111110000010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111110100110111100010100101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111110100111101001110101101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110001111100011001001011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110101011111101110110100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110111110001100010010110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111011011100101101110100100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111100001000110001110001011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111110000001101101010100110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111100100011000111010101011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111111000100010101011000001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b00111111000100101100001100010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111111000100101110010111010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b10111101101110101100000011010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111111000000001010001101111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111101100101101101010001011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111101011001110010100110111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b00111101100110110010010110000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111110110100110111000011001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111101010100000110010101110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111101101110101111011000100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b00111101100110110000011011100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111110101111001100010000001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111110110011101110111000010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111110100111011100110110111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111111001001000110111001010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111110001111001010000100110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111101011000001010111110001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b10111100100111111011001110100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111110111010011111000100011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b00111101110100000011011000100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111111000000010101010110001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b10111101010000101110101011111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111110110011101011110100100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111110101100101110111011100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b10111100000010010000000000001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b10111110011001001110100000010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b00111110000000100100111001110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b10111101001110110010100110010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111011111100000111111001101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b10111110011001101111010001101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b10111100000101100000111010000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel27_Valid_Out)
	);
	Adder_64input add_k27(
		.Data1(Data_Out_Kernel27[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel27[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel27[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel27[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel27[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel27[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel27[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel27[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel27[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel27[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel27[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel27[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel27[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel27[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel27[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel27[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel27[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel27[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel27[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel27[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel27[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel27[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel27[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel27[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel27[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel27[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel27[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel27[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel27[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel27[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel27[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel27[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel27[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel27[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel27[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel27[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel27[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel27[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel27[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel27[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel27[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel27[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel27[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel27[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel27[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel27[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel27[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel27[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel27[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel27[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel27[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel27[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel27[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel27[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel27[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel27[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel27[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel27[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel27[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel27[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel27[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel27[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel27[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel27[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel27),
		.Data_Out(add_k27_Data_Out),
		.Valid_Out(add_kernel27_Valid_Out)
	);
	Batch_Norm bn_kernel27(
		.Data_A(32'b00111110001100101110111111001001),
		.Data_B(32'b10111100101011101011000011010101),
		.Data_In(add_k27_Data_Out),
		.Valid_In(add_kernel27_Valid_Out),
		.Data_Out(bn27_Data_Out),
		.Valid_Out(bn27_Valid_Out)
	);
	Relu_Core rl_kernel27(
		.Data_In(bn27_Data_Out),
		.Valid_In(bn27_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(rl27_Valid_Out)
	);
//////////KERNEL28//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111101001101101010000000111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110001101000011011101101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110011100000111101011010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110010011001111001000000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111110011101110011010011100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110000010001001001110101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111111001011100100011000010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111101100100010100001110010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110110101001000100011111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111011110011101011010000101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111110100001000000101001111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111110111000011011100111011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110011010001011001011101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111110010011001010000010000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111101010010000010111010000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111110100000000111010111101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110110011100100001101001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111110000010010111100001110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111110001011111110001011101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111101010110111010000011001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111111000000000010111110001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111110010001101111001101000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111111000000010101001000011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111111001110110001100101001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111110100111100100101010100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111101110110000100110110000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110100101111010001111000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110101111110110001011111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111100100000001110000100111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111101111111100101001101110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111110111010000101110110000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111101111000100011101111010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111111010001101011110100010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b00111110111010110110111101101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111111000001101100110000111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111101101111110110110110001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111111001110101010101101000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111110010000101110111110100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b00111101110011111110001010000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111101001111001100111011111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111111000100110101001101011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b10111101010000110110110001001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111101000101000001111011110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b00111101111100010101111101111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111111000111011011011000010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111111000100001010001110101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111110001101100000001011011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111101001001100110001100000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111110101101111101001110111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111101111011101010101000100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111110000111011000011011111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111110101111101011111000011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b00111100111110111011000101101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111111001101111101000011011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b10111100001001100011110011110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111110111111010000110100111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111110100000001111010010010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111110001111110110001000110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b10111110010001101100100001100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b00111101101100011100010110101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111101100101111010010101011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b10111110110100101110000001000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b10111101011100000010110011111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111110100011001000101101110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel28_Valid_Out)
	);
	Adder_64input add_k28(
		.Data1(Data_Out_Kernel28[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel28[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel28[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel28[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel28[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel28[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel28[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel28[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel28[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel28[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel28[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel28[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel28[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel28[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel28[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel28[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel28[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel28[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel28[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel28[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel28[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel28[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel28[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel28[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel28[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel28[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel28[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel28[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel28[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel28[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel28[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel28[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel28[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel28[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel28[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel28[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel28[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel28[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel28[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel28[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel28[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel28[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel28[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel28[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel28[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel28[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel28[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel28[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel28[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel28[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel28[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel28[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel28[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel28[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel28[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel28[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel28[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel28[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel28[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel28[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel28[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel28[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel28[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel28[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel28),
		.Data_Out(add_k28_Data_Out),
		.Valid_Out(add_kernel28_Valid_Out)
	);
	Batch_Norm bn_kernel28(
		.Data_A(32'b00111110000000011000101001100100),
		.Data_B(32'b00111110011010111010101010110111),
		.Data_In(add_k28_Data_Out),
		.Valid_In(add_kernel28_Valid_Out),
		.Data_Out(bn28_Data_Out),
		.Valid_Out(bn28_Valid_Out)
	);
	Relu_Core rl_kernel28(
		.Data_In(bn28_Data_Out),
		.Valid_In(bn28_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(rl28_Valid_Out)
	);
//////////KERNEL29//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110100110111111100001011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111110100010011111011101100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110001011100011011101101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111111000000100001110100100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111101101001011001101111011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111010000011010111101010001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111100100110011010011010101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111101011000001010000001110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111110101101111001111111011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111101101000100011010100101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111101100011101110001110100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111101101011111001010010000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111101000010111011001001000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111110011100110101110101001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110000110010110111110010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111100010010111010100001010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111111100000010011100000110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110101000011010110100110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111110010110000111001000001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111101110100000000111011101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110001010001101101010001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111100100110111110110110011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111110010100001000010001111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111110110001010100000011001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111110100010010110000010111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111110100111111100011110111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111101000001101111100000010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111101010001001110110110110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111110010001001111011010111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111100110111101001110111100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111101011100110010011101001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111110110111100001101110111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b00111110010100101011110000000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b00111101111011001111011001100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111110101100110101101000011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b10111101100101110101101111101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b10111110110010111001110010101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111101111000111010001110001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111111000000101100001001100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b00111110010101011011101100010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b10111110111101001101011001001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b10111101110101000111011011100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111101011110011001111010110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111100011010000010001011101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b00111110101010000010010011001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b10111110101011010101001110111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b10111101111000000111001101011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b00111110010100011010000010101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111110100101111010000100010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111101111111110111101110111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b10111101101000010110010100101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b10111110110110001111111001000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111110010001000111001011011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b00111101111010011100010101110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111110010110100000001110011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b00111101001111001001110001010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b10111111000000111010100110100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b10111110011001101100100010010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b10111101101001101110100000011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111101100011101000011010010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b10111101100110000100111010101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b10111100100110011110001101101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b10111010101110111010010111110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111101111101100001110111101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel29_Valid_Out)
	);
	Adder_64input add_k29(
		.Data1(Data_Out_Kernel29[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel29[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel29[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel29[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel29[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel29[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel29[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel29[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel29[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel29[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel29[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel29[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel29[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel29[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel29[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel29[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel29[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel29[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel29[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel29[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel29[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel29[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel29[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel29[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel29[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel29[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel29[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel29[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel29[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel29[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel29[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel29[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel29[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel29[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel29[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel29[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel29[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel29[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel29[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel29[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel29[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel29[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel29[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel29[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel29[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel29[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel29[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel29[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel29[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel29[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel29[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel29[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel29[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel29[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel29[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel29[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel29[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel29[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel29[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel29[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel29[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel29[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel29[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel29[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel29),
		.Data_Out(add_k29_Data_Out),
		.Valid_Out(add_kernel29_Valid_Out)
	);
	Batch_Norm bn_kernel29(
		.Data_A(32'b00111110001100110110110000000110),
		.Data_B(32'b00111111100001100000111010110010),
		.Data_In(add_k29_Data_Out),
		.Valid_In(add_kernel29_Valid_Out),
		.Data_Out(bn29_Data_Out),
		.Valid_Out(bn29_Valid_Out)
	);
	Relu_Core rl_kernel29(
		.Data_In(bn29_Data_Out),
		.Valid_In(bn29_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(rl29_Valid_Out)
	);
//////////KERNEL30//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111101100101010110110111000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111101110011010110010101111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111101111011110011000111011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110110000001010111010011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111101111111101110010111100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111011100000101101110010100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111101110001111011101100110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111100100010010100000001011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111110111011000111111000011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111110001110011000000000101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111101001101111000110111010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111101100000001000011010110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111110010001110000000101010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111110001010110100110000001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110010100000010100000001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111101111001111001100011001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111111000010100001111010001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110010010011111011110101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111101010111101101111010101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111101111100101101100101111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110110100100100101011011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111101111011100001111011000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111101100001111101001110010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111110011101111111101011101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111110101100101101100110100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111110100011001011101011000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111101100011001110111100101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110000011001110110101010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111011010000011100000110000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111110101010111110110110101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111101101111111101011011111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111110100100100010110000101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b00111111000001110110011001111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111110010010101110011001100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111101001101100000111100110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b10111110010100011101001011101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b10111111010101100111000000110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111101101001111101100000000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111110110011101011111001011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b00111110010000101100101011010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b10111111000010011101111010110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b10111110110001010001001011011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b00111100110010000000100111101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b00111100111000100110111111011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b00111110110001110001100010111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111110000000000010100110010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b10111101011111000110001011001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b00111101010110111110101110000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111011110010100010010101101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111110011010110000000011110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b10111101010000110010001011010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b10111110011110101111010101011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111110010111101001011110100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b00111110100110000111101100011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111100110100110111101000010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111110010011110110111101101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b10111110010010000110111010110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b10111110010000111101110100110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111101111001011001001011011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111110000101111101000000011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b10111110001111101000100101111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111101110110110100111110111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b10111110010000110101010010111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b10111101100110001100010011111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel30_Valid_Out)
	);
	Adder_64input add_k30(
		.Data1(Data_Out_Kernel30[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel30[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel30[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel30[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel30[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel30[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel30[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel30[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel30[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel30[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel30[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel30[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel30[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel30[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel30[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel30[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel30[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel30[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel30[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel30[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel30[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel30[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel30[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel30[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel30[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel30[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel30[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel30[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel30[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel30[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel30[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel30[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel30[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel30[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel30[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel30[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel30[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel30[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel30[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel30[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel30[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel30[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel30[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel30[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel30[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel30[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel30[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel30[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel30[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel30[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel30[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel30[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel30[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel30[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel30[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel30[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel30[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel30[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel30[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel30[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel30[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel30[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel30[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel30[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel30),
		.Data_Out(add_k30_Data_Out),
		.Valid_Out(add_kernel30_Valid_Out)
	);
	Batch_Norm bn_kernel30(
		.Data_A(32'b00111110001101100100111101110100),
		.Data_B(32'b00111111000100001001000110110100),
		.Data_In(add_k30_Data_Out),
		.Valid_In(add_kernel30_Valid_Out),
		.Data_Out(bn30_Data_Out),
		.Valid_Out(bn30_Valid_Out)
	);
	Relu_Core rl_kernel30(
		.Data_In(bn30_Data_Out),
		.Valid_In(bn30_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(rl30_Valid_Out)
	);
//////////KERNEL31//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111110101110101100001010011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111101101010010111111010000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111101011000000000110111000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111101111011001111011110110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111101101101010100110010010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111101101000011001010010010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111110000011000101001011001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111110000110101001000000111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111101101100000010100010101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111110000000110101010111111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111101100010100100101110101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111101100111000110101111111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111100111111100001100010111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111100110010000110111000000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111101110110111001010001101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111110001001111111110000011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110101000111011101010101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111010111101010011001001000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110000110000000010011000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111011010110100100001000100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110011010011000100111100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111101101101000001011011110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110010000101000111011101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111110001100111100001101001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111101101101000101001111010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110100100000000011101000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110111101101111101001101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111101101111010110110001011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111110010001110001001000111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111101111110011100001010001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111110110101100100000101011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110100110000100000001001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111101100111101001000000110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b00111110100101101011110001011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111110101100010001111010001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b10111101000110110001111110010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111110011010011110000000101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111110000111011100011111100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b00111110001000110110101010000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111101110010011110011011000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111111000110010011001110101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111101111111101010111000000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111011000001101011111111111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111101100000110100100100111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111110010000100011000001110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111110110010111111111001100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111110010011001100010100111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111110001110011110001110101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b00111100000101001000010100111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b00111101101011000111110101000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111101101100101101010001001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111110000111110011110110111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b00111110011000100011101100010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111110111100100001011100000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111101101110101000011111100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111110011011101010101111001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111110110011111100001111001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111110000100101101000110101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b10111110010111111111111110000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b00111101110111011101101011110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111110000000101001101111100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111101011100001111010110001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111110101011101011111110001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111100101011000001001110101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel31_Valid_Out)
	);
	Adder_64input add_k31(
		.Data1(Data_Out_Kernel31[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel31[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel31[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel31[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel31[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel31[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel31[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel31[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel31[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel31[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel31[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel31[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel31[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel31[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel31[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel31[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel31[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel31[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel31[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel31[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel31[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel31[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel31[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel31[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel31[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel31[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel31[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel31[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel31[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel31[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel31[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel31[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel31[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel31[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel31[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel31[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel31[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel31[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel31[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel31[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel31[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel31[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel31[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel31[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel31[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel31[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel31[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel31[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel31[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel31[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel31[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel31[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel31[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel31[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel31[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel31[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel31[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel31[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel31[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel31[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel31[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel31[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel31[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel31[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel31),
		.Data_Out(add_k31_Data_Out),
		.Valid_Out(add_kernel31_Valid_Out)
	);
	Batch_Norm bn_kernel31(
		.Data_A(32'b00111110010111001001011100110011),
		.Data_B(32'b10111111001001000001011111001000),
		.Data_In(add_k31_Data_Out),
		.Valid_In(add_kernel31_Valid_Out),
		.Data_Out(bn31_Data_Out),
		.Valid_Out(bn31_Valid_Out)
	);
	Relu_Core rl_kernel31(
		.Data_In(bn31_Data_Out),
		.Valid_In(bn31_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(rl31_Valid_Out)
	);
//////////KERNEL32//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111101110000100110000011110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111011010011100101101101010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111101011001110100010010110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110010001101011111111110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111100011011101010110010011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111110010100010010100001110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111111000010110000111001010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111110000100111010001111000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110011110111010011010101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110001100000001011111111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111110011110001001100110000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110000101101100000001000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110100010011001001111110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111110100110010101000110101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111101000001111000101011010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111110010100011010100010000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111110101011011010110000101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110110001000010001101110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111111010001110010001011111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110001111011110111001010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110011010101011011101001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111110001000111100111100010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111101111110111100001101100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111101101011010011001101111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111110101111100101001101001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111110100100100000101011011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111110001001010110000010101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111101110001010100000101111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111101000001010110001011000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111111000011101110110100110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111100110000101111010110101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111111100101010101010001010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111101111111011111010001011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111110100100111011110100001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111111001010000100110101001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b10111101011101100000011011101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b10111111010000011010101101000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111111001011010001101010110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111111011011011100101110100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b00111110100111100011100010011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b10111110101110110111111001111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b10111110110100111101110110100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b00111011100010100101010001000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111110000010100001110100010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b00111110101000000101000110111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b10111101010010111100101011000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111110100001011010001111001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b00111110100001010111101111111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b00111110100011010110110100011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111110100000000100001100000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b10111110001110110011101001000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b10111110011111010100011001011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111110111001111111001111110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b00111101001001100100100010100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111110111001000100000010011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b00111100011100000000010011110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b10111110010001111111000110101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111110000000011011000000001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b10111110010110111001101111101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b00111111001001000101000001100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b10111110100000110110100110001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b10111100011111111110000111111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b10111110100001000110001000001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111110000000110110001110011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel32_Valid_Out)
	);
	Adder_64input add_k32(
		.Data1(Data_Out_Kernel32[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel32[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel32[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel32[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel32[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel32[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel32[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel32[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel32[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel32[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel32[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel32[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel32[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel32[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel32[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel32[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel32[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel32[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel32[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel32[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel32[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel32[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel32[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel32[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel32[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel32[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel32[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel32[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel32[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel32[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel32[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel32[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel32[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel32[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel32[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel32[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel32[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel32[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel32[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel32[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel32[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel32[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel32[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel32[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel32[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel32[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel32[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel32[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel32[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel32[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel32[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel32[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel32[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel32[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel32[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel32[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel32[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel32[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel32[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel32[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel32[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel32[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel32[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel32[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel32),
		.Data_Out(add_k32_Data_Out),
		.Valid_Out(add_kernel32_Valid_Out)
	);
	Batch_Norm bn_kernel32(
		.Data_A(32'b00111110000101110001011011011101),
		.Data_B(32'b00111111011011101111101011011010),
		.Data_In(add_k32_Data_Out),
		.Valid_In(add_kernel32_Valid_Out),
		.Data_Out(bn32_Data_Out),
		.Valid_Out(bn32_Valid_Out)
	);
	Relu_Core rl_kernel32(
		.Data_In(bn32_Data_Out),
		.Valid_In(bn32_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(rl32_Valid_Out)
	);
//////////KERNEL33//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111110100110110111111001010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111101010111010011011101000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110001111001010100100001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110110101111111110111010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111101100110000011101010110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110100000100111000010110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111110110100000010001011000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111011100110111011001110001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110100000001110100110011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110100011101001001111100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111110011110101001110000011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111100001110100110101100110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110000001110101110111000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111101111100100111000011110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110000011010101000011011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111110001101110010111001000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110010111100111111110001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110000011001011100010101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110100001000110111111111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111110000111001000110101100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111111000101011000100010111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111101111001001001100111110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111111001000001000100110011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111111000001110000111101011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111111001100001011010011101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110101010000101100111000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110100001111000010100001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111101101111011110101011111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111111000011011010000001101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111110100101011110110110011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111101001000111000110010110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110101011100100001101010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111111000010010111100101100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111101010010111101101000111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111110001100001000011011111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111110001010101101110110011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111111001001000111010000001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b00111110000001011110110010100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b00111111001101001111000001110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111110011011011101111100100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111111011010001011011000111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111110010110101011111011110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111110011010000101000001010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b00111111000011011011001110110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111110111011001011100010110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111110100010000100010111000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b10111101101010011000010111001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111101011110111011010101111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111110100111101110010110010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111101111111111001110011010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111110110010111100100111001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111100101011000110111111100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111101101110001101001101101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111111001101100100000011001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b10111100010111001100101001010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b00111101000110010101010011110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111110010111110010010010101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111110111010101110000010111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111100011110010011111101010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111110011100110110011100011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111110101110011010111001110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b10111110011000110000111101001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111110110111101001010101010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b10111110101101101110001110010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel33_Valid_Out)
	);
	Adder_64input add_k33(
		.Data1(Data_Out_Kernel33[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel33[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel33[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel33[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel33[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel33[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel33[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel33[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel33[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel33[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel33[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel33[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel33[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel33[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel33[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel33[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel33[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel33[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel33[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel33[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel33[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel33[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel33[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel33[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel33[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel33[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel33[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel33[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel33[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel33[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel33[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel33[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel33[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel33[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel33[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel33[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel33[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel33[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel33[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel33[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel33[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel33[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel33[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel33[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel33[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel33[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel33[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel33[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel33[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel33[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel33[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel33[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel33[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel33[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel33[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel33[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel33[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel33[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel33[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel33[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel33[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel33[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel33[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel33[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel33),
		.Data_Out(add_k33_Data_Out),
		.Valid_Out(add_kernel33_Valid_Out)
	);
	Batch_Norm bn_kernel33(
		.Data_A(32'b00111101111100100000010000001001),
		.Data_B(32'b10111110010011110001000000010010),
		.Data_In(add_k33_Data_Out),
		.Valid_In(add_kernel33_Valid_Out),
		.Data_Out(bn33_Data_Out),
		.Valid_Out(bn33_Valid_Out)
	);
	Relu_Core rl_kernel33(
		.Data_In(bn33_Data_Out),
		.Valid_In(bn33_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(rl33_Valid_Out)
	);
//////////KERNEL34//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111110000011010000110001100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110100101011000011101110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110010000000001111110101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110010111101100101101011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111011101010011010110010110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110100001111000100101000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111110111101011110111001011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111101100101110010000101110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111101110000100000010100111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111110000100010100100001001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110110000011001000101001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111101101101010010101111001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110100101001111001100101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111101101000101000110011001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111101001100110001111010100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111011100001111010011000000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110110111111100110101100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111110001110001110001000100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111110110010100000000010111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110101110010010101000010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111111000100011000011111101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111110100111011010110010000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111111000000001111101000101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111110011111001110111100100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111101011100000010100011110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110011111100100001001111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111111000100001001110101101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110101011011000100101001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111100110010010110011001010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111110010101101011111000001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111110100000000111111101001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110110010101001000000111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111111001011010000011101000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b00111110110101101001001110000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111111001001000110001101001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111100001000001000101100111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111110110111110001110100011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b00111100001101010110101000000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b00111110000001010101010111110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111101101011010001000101110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111111000011100111011000000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111110101001011100111000111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111100110001100110100111110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b00111101100001000111111101000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111111000110001101001101010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111110101001111011011011111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111111000010000111010101011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111110101001101101111000110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111110100000100110011001011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b00111110101011001110101101100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111110101001000111001010101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111110110111010111110011001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b00111110010000010101001010100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111110101001111000111010000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b10111100010111111011100010011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111110100101000111110010100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111101111010111010001010011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111101110011010000011100111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b10111101100000111001001000001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111101100111001101101001101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111110100100110001100111000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b10111110000111101101101011001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111110010111001010111100110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b10111101001001111110011001000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel34_Valid_Out)
	);
	Adder_64input add_k34(
		.Data1(Data_Out_Kernel34[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel34[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel34[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel34[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel34[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel34[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel34[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel34[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel34[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel34[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel34[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel34[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel34[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel34[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel34[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel34[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel34[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel34[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel34[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel34[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel34[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel34[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel34[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel34[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel34[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel34[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel34[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel34[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel34[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel34[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel34[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel34[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel34[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel34[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel34[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel34[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel34[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel34[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel34[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel34[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel34[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel34[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel34[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel34[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel34[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel34[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel34[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel34[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel34[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel34[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel34[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel34[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel34[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel34[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel34[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel34[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel34[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel34[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel34[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel34[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel34[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel34[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel34[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel34[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel34),
		.Data_Out(add_k34_Data_Out),
		.Valid_Out(add_kernel34_Valid_Out)
	);
	Batch_Norm bn_kernel34(
		.Data_A(32'b00111110000111010000001110000110),
		.Data_B(32'b10111111000010010100100000110110),
		.Data_In(add_k34_Data_Out),
		.Valid_In(add_kernel34_Valid_Out),
		.Data_Out(bn34_Data_Out),
		.Valid_Out(bn34_Valid_Out)
	);
	Relu_Core rl_kernel34(
		.Data_In(bn34_Data_Out),
		.Valid_In(bn34_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(rl34_Valid_Out)
	);
//////////KERNEL35//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111110110000110110110100011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111101001110000001010010101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110110010110001110010010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110100101001110011101111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111110000010011010110101111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111101101000001001110101000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111101110110111000111011011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111101010111000110001010111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111101111101101011010111111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111110011001010011001111000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111101000001001110111001011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111100110100001111100000001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111101011110010001111111100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111110100110110010010111000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110000101000111111001101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111101110000011010111000101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111101001010100010000000100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111011111101010000011111101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111101011010001110011111011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110011101010010100100101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110101001110100001101011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111010110001011111110101111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110100011001001011100010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111101111100110010010101010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111101100111111001001110101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110001111011101010100000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110110001100011110011111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111111000011011110101100000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111110010010001000000010100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111110100000001100010100010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111110001110011111011100000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111011101101010010010111101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111110111101000010101011100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b00111110110001000010101011010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111111001101001100001000010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b10111110011010110011000000100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111110100010000100011011101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111110001100000001110001010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b00111100010001110000000011000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b00111101101111111000110100010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111110111100100000100000001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111110010010110100100001111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b00111101011000000100011110110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111101001011001101000101000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111110100100011000000010001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111110100111100111011110010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111101010010000100111111000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111111000001111110001001100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111100101101010111110111110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111110000011111110101101100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111101011101110010011001110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111110110011010011110001111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b00111110100011101010010010111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111111000001111010011011110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111110010100101100110010111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111110110001011001000110010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111110101010001110100101111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111110001001000001011000110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b10111101111111011111110001010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b00111110001000101011100001101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111101101111001101111110100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b10111110001101011100101011010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b10111011100101110100111101101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b10111101011001110111101010001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel35_Valid_Out)
	);
	Adder_64input add_k35(
		.Data1(Data_Out_Kernel35[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel35[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel35[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel35[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel35[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel35[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel35[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel35[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel35[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel35[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel35[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel35[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel35[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel35[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel35[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel35[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel35[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel35[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel35[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel35[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel35[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel35[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel35[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel35[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel35[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel35[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel35[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel35[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel35[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel35[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel35[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel35[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel35[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel35[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel35[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel35[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel35[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel35[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel35[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel35[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel35[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel35[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel35[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel35[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel35[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel35[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel35[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel35[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel35[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel35[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel35[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel35[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel35[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel35[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel35[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel35[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel35[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel35[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel35[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel35[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel35[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel35[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel35[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel35[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel35),
		.Data_Out(add_k35_Data_Out),
		.Valid_Out(add_kernel35_Valid_Out)
	);
	Batch_Norm bn_kernel35(
		.Data_A(32'b00111110010110100101101010100110),
		.Data_B(32'b10111110101001100111000001111011),
		.Data_In(add_k35_Data_Out),
		.Valid_In(add_kernel35_Valid_Out),
		.Data_Out(bn35_Data_Out),
		.Valid_Out(bn35_Valid_Out)
	);
	Relu_Core rl_kernel35(
		.Data_In(bn35_Data_Out),
		.Valid_In(bn35_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(rl35_Valid_Out)
	);
//////////KERNEL36//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111101100110101010111010100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110010101111010100011101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111101010110100010000110010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110100100001000011011010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111110011000001001111011101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111101001111011101110010110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111110100011010011000011100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111101010000101100101101001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111111000001101100111010110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111110010011001110000111110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111111001110000010110000101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111001100101011111101101110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111110010001000100100010100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111110101010110111010110101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110001000000000011111000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111110000011111111001000010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110100100111101111110011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111101100101010000110110100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111111010100111000010111111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111101111010111101110001010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111111001000100100111101010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111110100011100000001110011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111100101000111010000110101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111110110001001000110111111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111110100111110001010011101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110111001000011111010110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111111000100100111011100101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111110000011001100000001100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111111000101001000001110100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110110001000000101111010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111110011110110011010000100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111111100011100001001111110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b00111101111101100001110010100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b00111110100001101010111100110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111110110100101111100011010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b10111100100101111101100011100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111110100111111111111101011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111011001010011100011110000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b00111110100100011001010100011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111110100001000010101011111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111111010001100111100101110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111110110100011001101101010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111110100001011100011010101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111110100110001110100110110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111110111110000001101001111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111100010000010110111101011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b10111110000001100011011011011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111110101111000101100111011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b00111101110000100101110000000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b00111110111001000110101111001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b10111110000011111111011101011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111110001111111000111000011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b00111110100010000000101000101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111110101010001101010011000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b10111101000111110000011100000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111110010110010111100001011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b10111110110001111101110101101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b10111101101101110111101000001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111101001001011100011010000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111110100010101101101001101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b10111101111100101001101111001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111110101001110001101010000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111110101110101101011000110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b10111110110101110010101001101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel36_Valid_Out)
	);
	Adder_64input add_k36(
		.Data1(Data_Out_Kernel36[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel36[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel36[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel36[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel36[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel36[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel36[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel36[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel36[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel36[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel36[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel36[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel36[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel36[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel36[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel36[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel36[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel36[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel36[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel36[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel36[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel36[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel36[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel36[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel36[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel36[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel36[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel36[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel36[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel36[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel36[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel36[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel36[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel36[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel36[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel36[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel36[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel36[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel36[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel36[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel36[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel36[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel36[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel36[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel36[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel36[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel36[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel36[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel36[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel36[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel36[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel36[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel36[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel36[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel36[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel36[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel36[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel36[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel36[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel36[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel36[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel36[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel36[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel36[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel36),
		.Data_Out(add_k36_Data_Out),
		.Valid_Out(add_kernel36_Valid_Out)
	);
	Batch_Norm bn_kernel36(
		.Data_A(32'b00111110001011010001101101000001),
		.Data_B(32'b10111110101010101000110111011001),
		.Data_In(add_k36_Data_Out),
		.Valid_In(add_kernel36_Valid_Out),
		.Data_Out(bn36_Data_Out),
		.Valid_Out(bn36_Valid_Out)
	);
	Relu_Core rl_kernel36(
		.Data_In(bn36_Data_Out),
		.Valid_In(bn36_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(rl36_Valid_Out)
	);
//////////KERNEL37//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111111000110000101001110100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111101101110111001011001000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110001011111101101110110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111111000011001000011011110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111110001001100100001111010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111101100111111010110100110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111101001011100101011110010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111110000110011110001111010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111101111110000001001000000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111101101010111111111110111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111101001111111011111111111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111100110101111010000110101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110011100011010001110111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111101111011010001101101110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110001001010101100011000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111101010100110000010111011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110100100011110001110100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110100000011100001111011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110011110001001100101101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111101101000101010101001111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110101101110011100001100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111110001101110010110101001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111111001011010000101010111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111110100100111000011111100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111110101000011100111000110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110101011001101010001100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110011110101100111111101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111110000101001010011111001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111110010010101000101110000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111110111001111001010001111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111101011001101000110110111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110110101011000111100111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111110100011111101010001011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111101101011111111001100001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111110101110110011100010000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b10111101110110000111110101011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111110100110111001100100001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111101010000110101000101110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b00111110111100011000001110110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111110100000111001100011101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111111001000011111000001011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111110100100001001111011100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111110101001011010011101100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b00111110001000011101001000011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111111000100101000111101100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111110010001100001101001110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b10111101011101010110000010001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111110001011001101101000111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111110001011000111011000110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111101111110111001000110001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111111000010010110001110101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111110001000000111011011011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111101010110100001101111111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111110111011101010010000100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111110000100101111001100110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b00111100110011010101100001100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111110001110011001100101011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111110100000001111111011000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111110100100101001101101110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111110111010010110000001100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111110011001011111111101001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111110001110100101011101011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111110101111111010000111100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b10111110100110111100001111110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel37_Valid_Out)
	);
	Adder_64input add_k37(
		.Data1(Data_Out_Kernel37[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel37[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel37[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel37[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel37[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel37[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel37[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel37[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel37[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel37[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel37[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel37[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel37[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel37[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel37[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel37[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel37[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel37[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel37[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel37[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel37[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel37[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel37[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel37[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel37[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel37[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel37[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel37[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel37[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel37[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel37[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel37[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel37[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel37[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel37[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel37[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel37[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel37[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel37[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel37[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel37[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel37[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel37[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel37[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel37[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel37[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel37[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel37[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel37[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel37[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel37[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel37[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel37[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel37[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel37[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel37[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel37[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel37[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel37[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel37[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel37[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel37[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel37[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel37[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel37),
		.Data_Out(add_k37_Data_Out),
		.Valid_Out(add_kernel37_Valid_Out)
	);
	Batch_Norm bn_kernel37(
		.Data_A(32'b00111110001010001010100100011100),
		.Data_B(32'b10111110100110001111010111011000),
		.Data_In(add_k37_Data_Out),
		.Valid_In(add_kernel37_Valid_Out),
		.Data_Out(bn37_Data_Out),
		.Valid_Out(bn37_Valid_Out)
	);
	Relu_Core rl_kernel37(
		.Data_In(bn37_Data_Out),
		.Valid_In(bn37_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(rl37_Valid_Out)
	);
//////////KERNEL38//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110100110011111110000011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111110010011001101000101000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110010111000010011010011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110010100001101110010110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111101011110000101000000011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110011000000100110111011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111110010100100010111010110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111100100100101010111111001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111100000110101011111111011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111101101010011010011011010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111100010000100111010101111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110000101010001100010100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111101111001001011100011110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111101101110011000110101111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110110010100100111001010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111110110101011111111111011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111110111001100110101011110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111110010101010001100001101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111110001110100111000011111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111101010000000110001000001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110010101110001000111101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111110010101000101010011111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111100100000001000100000011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111110100111111100110010011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111101000101011011001000110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111110110100001000011011110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111111000000111111101111111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111110010000000100010111010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111110011010001001001011000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110101001100000110001101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111110001001011001101111110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111110101010111110000110111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111110000111001010111101101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111110100101011011101110100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111111001101100001101011100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111110000101100111101100100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b10111100100010010000100100001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b00111101111110101101101111000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111110010111010000011011001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b00111101101010000010101001110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b10111111000001101111001010101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111101101101111001011101001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b00111101111111101101011110010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b00111110010101101011011001011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b00111110100000110111111111101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b10111110001110001000101001100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b10111110001100111110010110111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b00111110101100101010011011100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b00111100110000000001011010011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b00111100010000110111001010000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111101110100110111000110001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b10111110011100011010101100010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111101111100111001010001110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b00111110010010000001001111001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111101110101000110101011001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111101000000101110011001010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b10111110111001001000100001101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b10111110010111001000011000101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111101111110001000000011111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111101101111011011001001110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111101100100001100011110101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111110000110001110010110001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b10111110000111011110100011100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111110011011010011011010011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel38_Valid_Out)
	);
	Adder_64input add_k38(
		.Data1(Data_Out_Kernel38[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel38[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel38[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel38[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel38[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel38[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel38[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel38[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel38[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel38[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel38[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel38[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel38[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel38[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel38[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel38[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel38[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel38[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel38[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel38[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel38[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel38[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel38[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel38[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel38[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel38[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel38[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel38[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel38[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel38[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel38[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel38[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel38[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel38[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel38[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel38[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel38[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel38[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel38[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel38[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel38[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel38[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel38[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel38[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel38[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel38[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel38[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel38[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel38[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel38[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel38[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel38[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel38[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel38[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel38[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel38[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel38[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel38[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel38[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel38[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel38[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel38[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel38[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel38[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel38),
		.Data_Out(add_k38_Data_Out),
		.Valid_Out(add_kernel38_Valid_Out)
	);
	Batch_Norm bn_kernel38(
		.Data_A(32'b00111110011000010110010011101001),
		.Data_B(32'b00111110100110010111110000001110),
		.Data_In(add_k38_Data_Out),
		.Valid_In(add_kernel38_Valid_Out),
		.Data_Out(bn38_Data_Out),
		.Valid_Out(bn38_Valid_Out)
	);
	Relu_Core rl_kernel38(
		.Data_In(bn38_Data_Out),
		.Valid_In(bn38_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(rl38_Valid_Out)
	);
//////////KERNEL39//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111110111111101000110101111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111110101000110011010001000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111101111110100010111110000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110100111011001111100010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111110101111010001110010101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111101011111010110100001011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111110100001111101111100010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111110011100000001111001000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111110111011001000010010000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111110100111000110111111011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111110010101110011011111101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110101100100000101001001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111101111111010011000100111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111101001010000011011011010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111101101011010111011111110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111110001100011010111001111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111110100110000110010101011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110110100011001111000011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110001110010110111001001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110111000111000111100100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111111010101010111110000111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111110111101010010111101011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111110100001110111100100110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111111000001110011000000100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111110001101111100011010101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111110111101000000010100101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111110010001101010100110111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111100110000010110111111100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111101111001101001010011111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111110100110100011110011101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111110100110010101101000100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111110110110011001110000111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b00111110111000111000010111000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111110001111100100111110011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111101110001100111010010000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b10111110100010111111000111101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b10111111001001111110111110110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b00111110100011101011000110000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111110111101111100101111111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111101110100100101110110111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b10111111011010010000100000001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b10111110101100100100100010001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111101010001001011010001000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b00111101001011011000001100011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b00111110101110000101111111011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111110000001111100101111001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111101110111110110101101000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111110000000101101111110110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b00111101011000110011000000011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111101010100100111010010101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111100111110100110100001001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111101100110001101001101001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b00111101111010110011000011010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b00111111010101011101011011101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111110011101010100111111101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b00111101101111100000100110001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111110111100001101101001010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111110000010111011000100010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b10111101101110000111101010011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b00111110101100110010100010001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111101100000100111111101101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111110101101011110000000100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b10111110101111100010100010111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111110100110010011110101111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel39_Valid_Out)
	);
	Adder_64input add_k39(
		.Data1(Data_Out_Kernel39[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel39[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel39[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel39[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel39[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel39[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel39[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel39[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel39[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel39[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel39[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel39[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel39[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel39[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel39[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel39[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel39[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel39[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel39[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel39[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel39[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel39[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel39[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel39[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel39[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel39[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel39[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel39[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel39[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel39[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel39[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel39[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel39[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel39[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel39[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel39[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel39[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel39[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel39[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel39[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel39[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel39[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel39[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel39[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel39[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel39[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel39[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel39[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel39[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel39[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel39[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel39[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel39[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel39[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel39[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel39[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel39[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel39[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel39[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel39[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel39[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel39[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel39[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel39[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel39),
		.Data_Out(add_k39_Data_Out),
		.Valid_Out(add_kernel39_Valid_Out)
	);
	Batch_Norm bn_kernel39(
		.Data_A(32'b00111110000100110111001111101110),
		.Data_B(32'b10111110110100111101110111010001),
		.Data_In(add_k39_Data_Out),
		.Valid_In(add_kernel39_Valid_Out),
		.Data_Out(bn39_Data_Out),
		.Valid_Out(bn39_Valid_Out)
	);
	Relu_Core rl_kernel39(
		.Data_In(bn39_Data_Out),
		.Valid_In(bn39_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(rl39_Valid_Out)
	);
//////////KERNEL40//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111110010100110110101100001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111100100000110101110001001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111111000110011011010000111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110000001000100010101000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111110001011010011101001010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110011010111000110000100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111111100011011001100111101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111110100111011100100000001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111101000111101101011011110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111110010011011110011000000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111110110001000001100101100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111110111011010001100100011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111101100000110110110001100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111110001111101100011101100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110100100111100101000001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111110110000100100110011011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111111000010110001000101011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111110110100011001111111111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111100010010010101110101111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110000101010011100011111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111100100011111001011011100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111110001010100111100101011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111111010000100000100110101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111110011100111000110101110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111111000011010011100101101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111101101011000101101101110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111110001011010111001001100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111101100011010000001110101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111110001101010011010100000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111101110110100101110110100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111110100100010000111000011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110101101100000011001011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111101011100010100101011001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b00111110100111011101011110000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111111001011111101110100010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b10111110001010001101110101100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111111000111100101101111100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b00111110100010001001110010001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b00111110001101100111000110011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111110000111110101100100101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b10111101100111011101000100001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b10111110110001011101011111000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111011110111010000001100111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b00111101111100110110111100101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111110100010110011011010111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111110101000010000000100110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111101111110100101100001100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111110000010111111111111000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111111000010000010001111011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111001101001111011000000100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111110000000010111110010000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111110100111111100110110010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b00111111000001001011010001111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111101011101100011000001111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b10111110100010111110010011000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111110100100001111010010011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111111001011110000011001010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111110000110001001111001110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b10111110000000001000101100001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b00111111000010000001001110011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b10111101010000100000110011001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b10111110100110101011111101001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b10111100100001001000110011100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111110100100011110001101011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel40_Valid_Out)
	);
	Adder_64input add_k40(
		.Data1(Data_Out_Kernel40[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel40[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel40[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel40[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel40[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel40[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel40[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel40[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel40[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel40[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel40[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel40[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel40[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel40[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel40[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel40[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel40[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel40[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel40[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel40[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel40[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel40[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel40[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel40[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel40[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel40[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel40[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel40[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel40[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel40[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel40[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel40[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel40[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel40[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel40[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel40[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel40[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel40[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel40[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel40[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel40[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel40[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel40[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel40[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel40[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel40[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel40[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel40[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel40[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel40[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel40[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel40[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel40[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel40[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel40[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel40[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel40[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel40[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel40[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel40[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel40[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel40[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel40[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel40[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel40),
		.Data_Out(add_k40_Data_Out),
		.Valid_Out(add_kernel40_Valid_Out)
	);
	Batch_Norm bn_kernel40(
		.Data_A(32'b00111110000110000101111101111111),
		.Data_B(32'b10111110010000110011000100001110),
		.Data_In(add_k40_Data_Out),
		.Valid_In(add_kernel40_Valid_Out),
		.Data_Out(bn40_Data_Out),
		.Valid_Out(bn40_Valid_Out)
	);
	Relu_Core rl_kernel40(
		.Data_In(bn40_Data_Out),
		.Valid_In(bn40_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(rl40_Valid_Out)
	);
//////////KERNEL41//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111110111010110101100000011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111101110110011100010000110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110000011000111011111000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110110110110101110001010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111100010001101100100011101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110010000011100011000101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111101001010010010100110001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111101100100011100010011100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111100011000100111100010000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111100010001010111110001010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110010011010011111100101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111101000101011010011110001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111101100010011101001111011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111101111000100001010111111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110100101000000111101101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111100100110111011000100000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111111000011010100001111101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110000111010010110101111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110011000100000010101100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110001101011101100011001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110100100101110011000110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111110010001001100011011001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110101111111001011111010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111110001111001101100000110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111110011000010010000100110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110100011100110110011010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110011000010110101010011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111110010101001010011100100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111110000011100110001000110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111110110110001111000100100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111101100111001001000101001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110110000110001111011111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111101010101111111001111111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b00111101100101100001000111110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111110110001110000100010100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b10111101111111100101110100001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111110101011101010101101011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b00111101000111110110100100011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b00111110110001000011110000010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111101111100111100110111111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111111001010100001001100011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111110101001100110100110001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111101111101110011001111000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b00111011100101100011000011000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111110101100111101101010000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111110010011010110111101000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111101011111010110100110100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111110010000111010011000001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111110001011011101101001011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111110000100111110111011111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111110100000111111100111001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111101000010110010010100111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b00111100100011011111110110101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111110101011101100111011000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111110000011001100010101000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111100110000011000111001101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111110101000011010011001100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111110010111100000111101010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111110001011001110101100100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111110000100001000110011000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111110010101011111110011011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111101101000001000011011101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111110100001001100101010110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b10111110000001111011000011111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel41_Valid_Out)
	);
	Adder_64input add_k41(
		.Data1(Data_Out_Kernel41[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel41[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel41[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel41[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel41[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel41[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel41[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel41[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel41[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel41[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel41[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel41[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel41[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel41[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel41[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel41[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel41[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel41[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel41[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel41[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel41[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel41[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel41[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel41[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel41[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel41[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel41[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel41[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel41[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel41[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel41[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel41[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel41[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel41[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel41[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel41[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel41[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel41[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel41[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel41[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel41[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel41[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel41[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel41[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel41[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel41[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel41[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel41[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel41[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel41[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel41[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel41[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel41[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel41[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel41[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel41[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel41[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel41[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel41[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel41[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel41[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel41[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel41[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel41[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel41),
		.Data_Out(add_k41_Data_Out),
		.Valid_Out(add_kernel41_Valid_Out)
	);
	Batch_Norm bn_kernel41(
		.Data_A(32'b00111110001110101010010111101110),
		.Data_B(32'b10111111010000111110110001100001),
		.Data_In(add_k41_Data_Out),
		.Valid_In(add_kernel41_Valid_Out),
		.Data_Out(bn41_Data_Out),
		.Valid_Out(bn41_Valid_Out)
	);
	Relu_Core rl_kernel41(
		.Data_In(bn41_Data_Out),
		.Valid_In(bn41_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(rl41_Valid_Out)
	);
//////////KERNEL42//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111110000101001110110101110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111101100100100101010101101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111111001011110100101000001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111111001010010011110101111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111101001110010111000100010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111110101000000100000110111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111111001101101110100000011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111110001010110010011101101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111101001111010010111101011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111101101000101100110001001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111101111010011111100111010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110010001010110011110110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110011101010010000000100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111111000111101000111111010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110110101111011110101010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111101101111110101000001001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111110010101101000000010101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110110111100010011110011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111100111100101000101100110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110000010100100110101011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111100110011001001101101011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111110100111111101110100001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111110101010100111111001100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111110111101111000011010101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111100110110001001100110100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111110101000100110101110110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110010010100100101001101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110010110110111110111000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111110110101001010000110011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111110100001010000111000000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111100110101101011101011001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111111011011001000011101010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111111010011110100010011011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b00111100101010000110000101001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111110100100000010100000010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111110001000011001100010101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b10111111001000001110111100101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111110100000101011000000000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111111000101010111100100101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b00111101011001100100100010001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b10111110011010011001111110101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111110011100000101111100010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b00111110011111001110100001101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b00111110100001011110111001000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111101000001101101001000100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b10111110101011100111111110110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111110101011100010010110111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b00111101001000100100110111011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b00111110001111001010001011011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b00111101100110101001100010110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111100010110010100011000111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111101010001110101111110000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111110110011010011011111011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111110100000100100111010010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111111000100000101101111101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b00111111001100101111001010100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b10111101011100101011110111100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111110100000011000011100111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b10111101100100110111000100101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b00111010100100100000100101000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b10111101101110111011001000100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b10111101010111101100100011100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b10111110101101110011101001000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111110111100100101010111000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel42_Valid_Out)
	);
	Adder_64input add_k42(
		.Data1(Data_Out_Kernel42[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel42[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel42[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel42[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel42[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel42[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel42[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel42[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel42[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel42[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel42[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel42[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel42[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel42[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel42[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel42[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel42[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel42[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel42[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel42[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel42[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel42[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel42[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel42[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel42[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel42[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel42[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel42[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel42[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel42[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel42[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel42[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel42[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel42[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel42[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel42[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel42[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel42[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel42[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel42[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel42[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel42[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel42[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel42[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel42[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel42[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel42[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel42[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel42[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel42[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel42[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel42[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel42[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel42[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel42[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel42[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel42[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel42[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel42[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel42[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel42[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel42[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel42[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel42[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel42),
		.Data_Out(add_k42_Data_Out),
		.Valid_Out(add_kernel42_Valid_Out)
	);
	Batch_Norm bn_kernel42(
		.Data_A(32'b00111110001100101011001001000110),
		.Data_B(32'b00111111000010001000100110101100),
		.Data_In(add_k42_Data_Out),
		.Valid_In(add_kernel42_Valid_Out),
		.Data_Out(bn42_Data_Out),
		.Valid_Out(bn42_Valid_Out)
	);
	Relu_Core rl_kernel42(
		.Data_In(bn42_Data_Out),
		.Valid_In(bn42_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(rl42_Valid_Out)
	);
//////////KERNEL43//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111110110001111111000001011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110001111010001111100110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110101110000010100000110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110011011110101010101000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111101100101111010000010111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111101111110100111010111101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111110010001100110100011000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111100100111111001110000010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110100101000100011000101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111100000001010101110101000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110000010000001010100001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111110001010111100000110001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110001010000111011011011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111110011001000001100001000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111101010010111011101011110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111101010011101111011100100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111101011101000001100101000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111100101101111011111010000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111110001101000001000111001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110001001100010101110010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110101110110100100001001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111101100111011101001001001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110111000100010100010110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111110100111011000010100111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111110100011011011001010101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110100000001110000100011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110110101111111101111000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111111001010011000001110010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111110000111110010011101101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111110001011100100110110000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111110011100010011110111010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111100111110010110011101110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111111010110111010011010000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b00111110101101110100011001101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111111010100011000110101010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b10111101110111101001100011100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111111000001110001011011000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111110100101010100010101110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111110000101001110111110011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111101000111111110011001101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111110111101010110111001010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111101110100001000000110100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111110001001001001110001101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111001101001011101110000101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111111000001111100011011001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111110110111000101111011110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111110011001001010010010100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111110100101000110101010101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111110010010011110111111100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111101110000000011000110100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111110010101100100001011111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111110110111000110111011100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b00111110000111000100110001100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111111000100000111111000000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111110011010101001001010100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111110101101100101011010001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111110100001100010011110111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111110001110100111110011110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b10111110010000111011011111101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b00111110000100100111010110101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111101111101111000110000010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b10111110000010110110101000011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b10111100010000011110100010100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111101101101001010001010000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel43_Valid_Out)
	);
	Adder_64input add_k43(
		.Data1(Data_Out_Kernel43[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel43[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel43[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel43[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel43[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel43[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel43[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel43[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel43[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel43[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel43[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel43[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel43[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel43[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel43[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel43[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel43[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel43[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel43[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel43[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel43[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel43[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel43[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel43[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel43[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel43[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel43[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel43[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel43[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel43[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel43[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel43[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel43[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel43[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel43[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel43[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel43[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel43[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel43[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel43[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel43[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel43[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel43[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel43[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel43[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel43[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel43[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel43[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel43[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel43[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel43[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel43[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel43[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel43[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel43[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel43[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel43[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel43[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel43[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel43[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel43[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel43[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel43[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel43[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel43),
		.Data_Out(add_k43_Data_Out),
		.Valid_Out(add_kernel43_Valid_Out)
	);
	Batch_Norm bn_kernel43(
		.Data_A(32'b00111110001011011011110010010001),
		.Data_B(32'b10111100101100000010110000010111),
		.Data_In(add_k43_Data_Out),
		.Valid_In(add_kernel43_Valid_Out),
		.Data_Out(bn43_Data_Out),
		.Valid_Out(bn43_Valid_Out)
	);
	Relu_Core rl_kernel43(
		.Data_In(bn43_Data_Out),
		.Valid_In(bn43_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(rl43_Valid_Out)
	);
//////////KERNEL44//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110110011101000100010110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110000110111010010101000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111111000011001100000100011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111101101100110010001101100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111110100101111010100110111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111101010000001100000110011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111111001100000110011111000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111111001111010100001100000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111110000100001001001000011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110101001000110001111010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110100110000111111100100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110111001111101100011001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111111000011100111110011000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111110000110010011111100010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111101000001000100010111001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111111001001011010101000101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111101011011101110001100000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110100100000000010111001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111101101100010101101101011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110101110001100000110001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110010010111010111000111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111110110110011000011100101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111010101010101101011100100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111110100000100111110111010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111111000110111111111000111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111111000100010110001001111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111101000100110101111010111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110011100001000100100011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111110100010000110010000101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110111111001100110011010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111101100000110100100100111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111100111100111010111100110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b00111100110011011111111011000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b00111101000110011100000100000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111110110000111111100011100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111110001111111100011000000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b10111110100111001011100010000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111110000101010111010000010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111110100001111101001100010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111101100001100001010100000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111110011111101110110000100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111110101111010111010000010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b00111110011100001111000111011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b00111110000110100110010101111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b00111100110001111111110101110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b10111111000001111011100110100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111101101000101000011001100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b00111110010111110101110101110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b00111110100111010001000110011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b00111110010000100011111111010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111110111001001010110111111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b10111110000001011110110000110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111110110001011001010001000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111101101110111101101011111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111110111110101000111001010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b00111111010100010000110010101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b10111111001001111100001101110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111110001100001101110011110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b10111110011000001010111100100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111110101100101110111111011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111110100110101000111111101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111110011000001001100100110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111110110011111100110110111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b10111110101010111010010111110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel44_Valid_Out)
	);
	Adder_64input add_k44(
		.Data1(Data_Out_Kernel44[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel44[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel44[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel44[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel44[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel44[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel44[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel44[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel44[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel44[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel44[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel44[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel44[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel44[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel44[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel44[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel44[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel44[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel44[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel44[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel44[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel44[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel44[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel44[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel44[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel44[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel44[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel44[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel44[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel44[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel44[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel44[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel44[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel44[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel44[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel44[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel44[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel44[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel44[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel44[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel44[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel44[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel44[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel44[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel44[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel44[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel44[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel44[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel44[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel44[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel44[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel44[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel44[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel44[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel44[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel44[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel44[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel44[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel44[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel44[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel44[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel44[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel44[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel44[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel44),
		.Data_Out(add_k44_Data_Out),
		.Valid_Out(add_kernel44_Valid_Out)
	);
	Batch_Norm bn_kernel44(
		.Data_A(32'b00111110010010001001100001111001),
		.Data_B(32'b10111111000101000000000011000111),
		.Data_In(add_k44_Data_Out),
		.Valid_In(add_kernel44_Valid_Out),
		.Data_Out(bn44_Data_Out),
		.Valid_Out(bn44_Valid_Out)
	);
	Relu_Core rl_kernel44(
		.Data_In(bn44_Data_Out),
		.Valid_In(bn44_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(rl44_Valid_Out)
	);
//////////KERNEL45//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111101111111110001110100111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110101111011010100100011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110000110010111000000010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110010110001101000010111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111110100100110101100111101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110010001110001000001000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111110111010010010011001101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111110000001111110001101010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111111001111001000110011100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111110011111100000101011101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110111000011111101110100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111101010001110100100000100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111101000000101110001110110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111101110000111000100111010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111101101010001010010100110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111110010000111011011101011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111111000101010001110110100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111110001000010011110011111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111111000010100100000010011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110101001110110101111100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110110111011110111101101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111110101101001100001000011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111101011110010111110111000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111111010101010101010101001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111101011100100111111011100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111110000000100001111001111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111111000001111100011101110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111101000000010001111101000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111111000011111100100111000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110100110110101100111010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111110100001011011001000111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110110101001010011011111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111110100000101010010000000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b00111111000111101110010011101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111110111001111111101101110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b10111101101100000011111011011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111110111110000101110010010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111101101100000111011000100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b00111110011011000011000110001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111101010011001000000001110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111111000110100101010101111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111101100001001100010101101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111101000011010100111010000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111110010111011010000000101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111110110000100000101101110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111110110111101001010111110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111110000010000100111001100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111111000010110111110100000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111110010110011100100000001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b00111110000110010000111001100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b10111110001001000101001000111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111110101011101100000100001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b00111110100001010101010111010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111110111011111011110101101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b10111110001000011110110011101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111111001011011010111110000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111011110110111001011010010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b10111110001000001001111001001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b10111110010010111111010000101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b00111110100011110011111011110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b10111011100110110110101111111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111110001000110101010110110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111110000001100101011100001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b10111101001011011111101111001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel45_Valid_Out)
	);
	Adder_64input add_k45(
		.Data1(Data_Out_Kernel45[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel45[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel45[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel45[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel45[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel45[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel45[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel45[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel45[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel45[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel45[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel45[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel45[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel45[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel45[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel45[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel45[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel45[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel45[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel45[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel45[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel45[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel45[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel45[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel45[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel45[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel45[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel45[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel45[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel45[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel45[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel45[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel45[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel45[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel45[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel45[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel45[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel45[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel45[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel45[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel45[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel45[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel45[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel45[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel45[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel45[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel45[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel45[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel45[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel45[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel45[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel45[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel45[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel45[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel45[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel45[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel45[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel45[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel45[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel45[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel45[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel45[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel45[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel45[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel45),
		.Data_Out(add_k45_Data_Out),
		.Valid_Out(add_kernel45_Valid_Out)
	);
	Batch_Norm bn_kernel45(
		.Data_A(32'b00111110000010110111111110000011),
		.Data_B(32'b10111110010101101100110000010101),
		.Data_In(add_k45_Data_Out),
		.Valid_In(add_kernel45_Valid_Out),
		.Data_Out(bn45_Data_Out),
		.Valid_Out(bn45_Valid_Out)
	);
	Relu_Core rl_kernel45(
		.Data_In(bn45_Data_Out),
		.Valid_In(bn45_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(rl45_Valid_Out)
	);
//////////KERNEL46//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110100001000010111000000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111111000111100110011010011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110101100110000011001010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110111010100000010111111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111110000111011111101101001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111101011111001001100110010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111110010100001100101001100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111101110000100110100111100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111101110001111010011110100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110000011110010001100001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111101101000011011111011010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111101010111101110000111101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111101011001100100100000100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111100111111110101011111000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110100101111011011110011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111101101101111011110000100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111111000001110111111011111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111101001010010100110000010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110100101101100011111011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110000000111001001001110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110100011001110100101001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111100110111010110001001011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111110111100011001011011001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111110100001010010111110000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111101010010010000010010010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111110010101110000111111011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111110011011101001011010110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111110101000000010101010101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111110011001011100101011110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110000011010011100010010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111110001011111011100110111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111111000010110000011000010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b00111101101111100000110000001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111110100100000110011101110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111110101001110110010011000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111110010001110110101100111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b10111110110010010110000110001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111101110110011101000000110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111110110000100000010000000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b00111101011110011000000101001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b10111111011001001100011000001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111101000010110110110100101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b00111110000100001110100111101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b00111100100011110011111000000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b00111110101010000011111100111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b10111110011100100111011011111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b10111110000101011010111010000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b00111110001100011010111011110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b00111101001010001011101000010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111101110010001010100101010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b10111011111001101111010010110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b10111110100101100100100011101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111110101101001001111101010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b00111101100100010000110001010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b10111100000110001010111111001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111101101010101000110001010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b10111110101000100110011001001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b10111110110001000110011110011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111101110010001111110010010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111110010010110000110001110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b10111110100110000101111101111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111100111001101110001000010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b10111110000011101000111001111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111101110111000010000001001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel46_Valid_Out)
	);
	Adder_64input add_k46(
		.Data1(Data_Out_Kernel46[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel46[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel46[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel46[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel46[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel46[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel46[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel46[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel46[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel46[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel46[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel46[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel46[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel46[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel46[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel46[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel46[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel46[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel46[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel46[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel46[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel46[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel46[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel46[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel46[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel46[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel46[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel46[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel46[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel46[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel46[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel46[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel46[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel46[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel46[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel46[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel46[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel46[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel46[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel46[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel46[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel46[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel46[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel46[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel46[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel46[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel46[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel46[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel46[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel46[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel46[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel46[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel46[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel46[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel46[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel46[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel46[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel46[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel46[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel46[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel46[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel46[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel46[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel46[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel46),
		.Data_Out(add_k46_Data_Out),
		.Valid_Out(add_kernel46_Valid_Out)
	);
	Batch_Norm bn_kernel46(
		.Data_A(32'b00111110001001001111101110000001),
		.Data_B(32'b00111111011101100001110000110100),
		.Data_In(add_k46_Data_Out),
		.Valid_In(add_kernel46_Valid_Out),
		.Data_Out(bn46_Data_Out),
		.Valid_Out(bn46_Valid_Out)
	);
	Relu_Core rl_kernel46(
		.Data_In(bn46_Data_Out),
		.Valid_In(bn46_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(rl46_Valid_Out)
	);
//////////KERNEL47//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111011111001011000111010110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110101100100000110101110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110000000010000100101011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110001000111010100110101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111110001111001000011011111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111011100101000100011100000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111110011010011101010011100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111110111100101010001010101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111101100111000000100010001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110010001011111001011110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111101100110010111010000001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110100101011010101011111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111111011010011110111000101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111110001110010000000011101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111101100110110000100101100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111111000010011110011000111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110001000100111101101000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111101001001111111000001100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110011100111111000010001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110001110001100000000100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110111111111111101000111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111110110111100011110011111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110110111000100110011111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111101100111101011101010010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111100101110101110010001010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111111000010000100101110111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111100100000101010001110110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110011101101010000111111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111111011010000101110000111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110011011110010100110011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111101110101000000111101111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110001001111010101111011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111111000000000010001011100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b00111101100101000101110110010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111110000110000101100000100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111110100100100010011110001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111110101000010111011011110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111110000000001100010111101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111101110100100111100101011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b00111110001111100001001100100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111110101010100100011000101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111110101001100001110101011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111101110010010011110001101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b00111110101101011111110100101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111110111010000011111000100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b10111100101100111010111111101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111110110110000111000011010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b00111110000010000100100010010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b00111101011000001100010011000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b00111110001101011011010001001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111111000111110001111011111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111101100110101111010111111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111110101110111100101100000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111110111001111000101100110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111110110111100111001110000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b00111111010000101100010000010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b10110101101100001110011110000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111110101111101101001111010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111110001101101001111101100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111110000001110101011011001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111111000011101001100110001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b10111110010111111000110101010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111110110111100000100011101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b10111110110000100010101011001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel47_Valid_Out)
	);
	Adder_64input add_k47(
		.Data1(Data_Out_Kernel47[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel47[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel47[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel47[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel47[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel47[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel47[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel47[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel47[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel47[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel47[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel47[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel47[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel47[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel47[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel47[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel47[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel47[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel47[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel47[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel47[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel47[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel47[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel47[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel47[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel47[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel47[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel47[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel47[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel47[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel47[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel47[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel47[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel47[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel47[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel47[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel47[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel47[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel47[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel47[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel47[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel47[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel47[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel47[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel47[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel47[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel47[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel47[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel47[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel47[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel47[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel47[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel47[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel47[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel47[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel47[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel47[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel47[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel47[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel47[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel47[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel47[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel47[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel47[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel47),
		.Data_Out(add_k47_Data_Out),
		.Valid_Out(add_kernel47_Valid_Out)
	);
	Batch_Norm bn_kernel47(
		.Data_A(32'b00111110011100011111010101010001),
		.Data_B(32'b10111111100011100110110000011100),
		.Data_In(add_k47_Data_Out),
		.Valid_In(add_kernel47_Valid_Out),
		.Data_Out(bn47_Data_Out),
		.Valid_Out(bn47_Valid_Out)
	);
	Relu_Core rl_kernel47(
		.Data_In(bn47_Data_Out),
		.Valid_In(bn47_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(rl47_Valid_Out)
	);
//////////KERNEL48//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111110010001100110101010011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110001110101000000000011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110100000011011101011010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110110111000001010001110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111100000011010000100010000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110100101000110101100100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111100011111110100101101101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111110110011001110010100000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111100001111101110001111110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111100100000101010001000110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111110001110001101011110001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111110000011001110111000010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110000100101111001000111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111101111010000011110100011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111111000101011001001010000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111101000100100101111110010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110001001001110011001100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111101001110010111101110101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110100110011110101111100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110111010111001011110011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110101001000101101110100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111101001010011101110111000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110101100001011110000100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111110011101110000100001111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111101011100010100010111011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111101111010110011011110110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111101110101001101100101011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110001101110110110010100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111110010000000010111000110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111111000101101101001110100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111110010001001110111001010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110001101100101100110111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111101001001011111010011101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b00111101111100111000011111011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111110100100000010101010001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b10111110001111100101100111010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b10111110000000100000000011110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b00111101110111011111011100110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b00111101011111100100111110110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b00111110010110011101011010000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111110111110100111100111010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111110010110000000000011010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111100100110010010100000010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111110001111000011100111010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111110100111010000010110110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111101110111001100000011101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111110000001011010110001001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111110110110011010100101110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111101100011110000011110011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b00111101000100001110010010001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111110110111001100100010011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111110010101001001010000000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b00111101000011101000001101010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111110100001011111111110110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b10111101110011111110101010001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111101001001000010111011001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111110001101101100101000110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b10111101010101000100000110011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111101100100010100000110100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111110010100101001111001011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111110010000011001000100101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b10111101000011001011001110010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111110000001111010111111010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b10111110001011101111101110011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel48_Valid_Out)
	);
	Adder_64input add_k48(
		.Data1(Data_Out_Kernel48[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel48[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel48[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel48[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel48[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel48[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel48[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel48[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel48[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel48[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel48[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel48[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel48[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel48[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel48[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel48[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel48[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel48[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel48[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel48[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel48[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel48[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel48[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel48[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel48[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel48[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel48[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel48[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel48[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel48[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel48[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel48[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel48[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel48[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel48[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel48[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel48[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel48[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel48[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel48[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel48[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel48[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel48[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel48[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel48[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel48[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel48[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel48[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel48[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel48[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel48[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel48[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel48[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel48[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel48[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel48[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel48[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel48[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel48[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel48[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel48[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel48[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel48[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel48[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel48),
		.Data_Out(add_k48_Data_Out),
		.Valid_Out(add_kernel48_Valid_Out)
	);
	Batch_Norm bn_kernel48(
		.Data_A(32'b00111110100010110011100110001010),
		.Data_B(32'b10111110010010011010010011110011),
		.Data_In(add_k48_Data_Out),
		.Valid_In(add_kernel48_Valid_Out),
		.Data_Out(bn48_Data_Out),
		.Valid_Out(bn48_Valid_Out)
	);
	Relu_Core rl_kernel48(
		.Data_In(bn48_Data_Out),
		.Valid_In(bn48_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(rl48_Valid_Out)
	);
//////////KERNEL49//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111110000100011101101100111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111101000101101010000000001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110101110110111011111000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110010011100001100110111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111110000011110010101010000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110111100110110100100001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111111000111100110110010110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111110010011101001111101011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110110000001111111001100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111110101100110010110100111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110101001111111101001101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111101111101110000101000000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111101101010101000111111000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111110100101101011000111001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110100001001111000110000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111110101010010110000101110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111111000011001100110101111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111110001100010110010011101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111110100010000100101111100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110001100111011000001011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110001001101011011110100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111110100011001111110101110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111111000000010011010000010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111111010001001110001010111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111110010000011011000010011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111011001010101110000001000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110100010011010100100101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111100110010100001001100101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111111001000110000111000110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111100001011001101111011110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111110010001111101101100110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110101100010000101011110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b00111110011001010110011110011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b00111110110111011010000110111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111111001011000110110110011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b10111110110101111111111000111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111110101010111010100101010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b00111100111101010100010000111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111101101010111110110001010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111110010011101000101000000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111100101100011000110101110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b10111110001100010010000100011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111110001001100111101000101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111010100010011010100111100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111110110011011101000001000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111110011110101100101111010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b10111100101011100110010000101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111110000111010001100101110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111110110101011001000001100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111110000011111010100111001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111110100011011110110001001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111101111100100000100110101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b00111111001011101001101011011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b00111110110111010110000110111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111110110110111001001111110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111111000001001011001010111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111111010000111111010011001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111101011101101010101110010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b10111110101100000110111001000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b00111111010111110000110111010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b10111101000111110001010111100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111101101011100000100001010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111110011101101000110011100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111011111010101010010010011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel49_Valid_Out)
	);
	Adder_64input add_k49(
		.Data1(Data_Out_Kernel49[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel49[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel49[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel49[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel49[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel49[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel49[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel49[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel49[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel49[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel49[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel49[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel49[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel49[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel49[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel49[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel49[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel49[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel49[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel49[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel49[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel49[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel49[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel49[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel49[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel49[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel49[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel49[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel49[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel49[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel49[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel49[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel49[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel49[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel49[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel49[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel49[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel49[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel49[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel49[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel49[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel49[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel49[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel49[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel49[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel49[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel49[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel49[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel49[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel49[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel49[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel49[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel49[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel49[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel49[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel49[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel49[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel49[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel49[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel49[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel49[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel49[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel49[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel49[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel49),
		.Data_Out(add_k49_Data_Out),
		.Valid_Out(add_kernel49_Valid_Out)
	);
	Batch_Norm bn_kernel49(
		.Data_A(32'b00111110000100111011011001011011),
		.Data_B(32'b10111110001111000010010100011100),
		.Data_In(add_k49_Data_Out),
		.Valid_In(add_kernel49_Valid_Out),
		.Data_Out(bn49_Data_Out),
		.Valid_Out(bn49_Valid_Out)
	);
	Relu_Core rl_kernel49(
		.Data_In(bn49_Data_Out),
		.Valid_In(bn49_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(rl49_Valid_Out)
	);
//////////KERNEL50//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110111010100001011001010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111101011010001010110011001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111101110010001000101011111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110100101011101011110111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111101110010011100001101001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110000101010101110011110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111110010111011010011001101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111110100110011101000110110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111111001010100001110101000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110011011010110100011111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111111000001010001010001011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111100110001111000001111100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111101111011010000001101001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111110100110100110110100011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110101101100111011110110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111111010101011001010111101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111110110110101000100010011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111101100101110100011001000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110001001001000011001011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111011110111100001000111010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110101111010101110001011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111110001110000100001101011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111110001110101001011111000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111111010100111111011101111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111110100000100110010100000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111101100010110001100110111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111110111000010001011001000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111111000010001011000001010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111101110111110110000101111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110011011000111101010101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111100100110011011010100110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111110010111011001000101110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b00111110100010101011010101101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111110010101101100111101000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111111001011000001100010110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b10111101001010000101110110110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111101001110110100101111000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111110001010010100001101001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111111000100101001101110110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b00111110100000000110110111011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b10111111000001110101001000011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b10111110100111001011001111110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b00111110000110101010001111110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111101111100001000010111010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b00111110101010000011011010000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b10111110111100101010000111101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111101110100001101100010100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b00111110110101111110001101110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b00111101110110010101111111110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111101100111010111101100000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111101110001010110101000111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b10111110101111011010011000001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111101101111010011111000101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b00111110111111100000101110011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b10111100001100101000100101011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b00111101101111000100100010111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b10111111000010010110100100100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b10111110011100010110100000001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b10111110001001100001000110110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b00111110001001111010001001010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111100001011100011100000001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b10111110101111000100100000101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b10111101001110101000000011001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111101000100101101011001101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel50_Valid_Out)
	);
	Adder_64input add_k50(
		.Data1(Data_Out_Kernel50[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel50[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel50[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel50[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel50[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel50[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel50[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel50[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel50[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel50[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel50[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel50[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel50[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel50[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel50[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel50[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel50[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel50[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel50[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel50[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel50[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel50[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel50[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel50[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel50[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel50[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel50[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel50[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel50[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel50[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel50[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel50[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel50[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel50[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel50[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel50[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel50[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel50[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel50[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel50[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel50[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel50[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel50[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel50[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel50[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel50[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel50[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel50[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel50[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel50[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel50[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel50[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel50[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel50[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel50[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel50[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel50[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel50[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel50[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel50[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel50[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel50[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel50[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel50[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel50),
		.Data_Out(add_k50_Data_Out),
		.Valid_Out(add_kernel50_Valid_Out)
	);
	Batch_Norm bn_kernel50(
		.Data_A(32'b00111110000010000100110010101010),
		.Data_B(32'b00111110111110101101111100001010),
		.Data_In(add_k50_Data_Out),
		.Valid_In(add_kernel50_Valid_Out),
		.Data_Out(bn50_Data_Out),
		.Valid_Out(bn50_Valid_Out)
	);
	Relu_Core rl_kernel50(
		.Data_In(bn50_Data_Out),
		.Valid_In(bn50_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(rl50_Valid_Out)
	);
//////////KERNEL51//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111100011111011110110100101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111110001110010110101100110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110110101110000101100100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111111000110001110001110010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111100111011011010000001101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111110110110111101110100010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111110100000010101001111100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111110011010000000000110110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111110000111111010000100011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111110100010000100111000101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110001110001000110110111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111101110011101010010111111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111101110100100101001010101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111100101110001101101000111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111101000110011001100000000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111110110110111111100011001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111111000010100111101000001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110100010011110110001000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111110010100100011110001110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111101100001000010001010100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110101011111110010001110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111110100011001110100011110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111111011001001101100110011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111111000001010010000100111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111110101001000001010000111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111111000101010010000101011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110100111010110101000100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111110101000111101100000101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111100001100101110100001110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111110001011000111000001111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111101111011001001011001100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111111000010011101111111111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111110100100010101110000001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111110010110010011010000001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111110101010010110000010100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111101010000000011101010100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b10111111011101101001000100010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111110011010010000001010001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111111000101100001011000001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b00111110011010011001110111010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b10111111001111101001011101001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b10111110000011011110110000100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b00111110100101111011010010010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111110011101000010110001000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b00111110101110001100100000011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b10111101010011111000000110100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111101101100000010100101001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b00111100100001010100011100011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b00111110010011100000110010001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b00111110010110111010111001111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b10111110101110001011101010100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111100001010011111111010111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111110100010101101001100111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b00111101100010001100011100110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111101001100110001100111000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111100011110100010111000100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b10111110000101100011101010100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b10111110000010101111101000100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111100110000000100011100111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111110100000011110100000011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b10111110101010110001011010010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b10111100101010111101101101000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b10111111011001101001000010100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111110110110001011111001011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel51_Valid_Out)
	);
	Adder_64input add_k51(
		.Data1(Data_Out_Kernel51[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel51[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel51[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel51[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel51[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel51[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel51[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel51[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel51[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel51[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel51[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel51[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel51[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel51[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel51[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel51[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel51[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel51[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel51[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel51[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel51[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel51[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel51[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel51[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel51[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel51[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel51[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel51[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel51[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel51[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel51[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel51[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel51[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel51[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel51[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel51[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel51[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel51[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel51[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel51[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel51[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel51[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel51[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel51[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel51[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel51[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel51[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel51[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel51[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel51[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel51[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel51[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel51[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel51[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel51[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel51[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel51[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel51[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel51[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel51[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel51[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel51[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel51[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel51[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel51),
		.Data_Out(add_k51_Data_Out),
		.Valid_Out(add_kernel51_Valid_Out)
	);
	Batch_Norm bn_kernel51(
		.Data_A(32'b00111110000000110001100001110001),
		.Data_B(32'b00111111011000111011000010111110),
		.Data_In(add_k51_Data_Out),
		.Valid_In(add_kernel51_Valid_Out),
		.Data_Out(bn51_Data_Out),
		.Valid_Out(bn51_Valid_Out)
	);
	Relu_Core rl_kernel51(
		.Data_In(bn51_Data_Out),
		.Valid_In(bn51_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(rl51_Valid_Out)
	);
//////////KERNEL52//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110110000111011111010111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111101110100100011100101011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111101110000001001101100100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110111011000101110100101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111101101011001100001100011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111101000111100111101001010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111110001111001011100011111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111110000110111100100011001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111111000010010011111000101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111101001001110010010101110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111101110101101101000011101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110010101101101101100011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111100111000110001001010100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111101101001101000111111000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110101100110010111110000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111100000001100011011110000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111111000011001100000100010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111100101001110100110000110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111110011010101010011110110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111101100101100010000111111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110100011111100011001111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111100100001100110111010100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111110100000111010001100101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111110001110000111111110110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111110010111101010111011101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111110100001110100111010111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111110000111010110010101011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111110100110100010001000010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111101100010111000001100000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110010101010101010100111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111101000100001011111110100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111110000101011001111011111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b00111110100110100100101001101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111110001011010000011111001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111110111110000110000011010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111101010101000110100001011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b10111110110000010010001100011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111101101000100011001101101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111110110010000110110111100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b00111101101001011011001100011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b10111110110010100111010000111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b10111101101111100010010000011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b00111110000011000010011111000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b00111100101100000001000100100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b00111110100101101110101101111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b10111100101111110011110010101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b10111101111101111000100100001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b00111110100101100101101010110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b00111101011001011010100000001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111100100011111111101000011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111110000101000110001001101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b10111110010111110110110010110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111101011010011001111011010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b00111110100000000001000110110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111101001110100010001011100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b00111100000110101100001011011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b10111110101001011000101011101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b10111110111010101010001001001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111110010100011100011100101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111110000000011001011011000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b10111101110111110010001001011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111101110110010011001000011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b10111100110001100110100101101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111110010100000000010111000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel52_Valid_Out)
	);
	Adder_64input add_k52(
		.Data1(Data_Out_Kernel52[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel52[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel52[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel52[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel52[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel52[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel52[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel52[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel52[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel52[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel52[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel52[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel52[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel52[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel52[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel52[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel52[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel52[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel52[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel52[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel52[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel52[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel52[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel52[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel52[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel52[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel52[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel52[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel52[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel52[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel52[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel52[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel52[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel52[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel52[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel52[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel52[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel52[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel52[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel52[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel52[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel52[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel52[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel52[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel52[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel52[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel52[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel52[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel52[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel52[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel52[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel52[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel52[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel52[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel52[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel52[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel52[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel52[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel52[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel52[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel52[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel52[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel52[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel52[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel52),
		.Data_Out(add_k52_Data_Out),
		.Valid_Out(add_kernel52_Valid_Out)
	);
	Batch_Norm bn_kernel52(
		.Data_A(32'b00111110010010010010101001001111),
		.Data_B(32'b00111101101001010110010101111000),
		.Data_In(add_k52_Data_Out),
		.Valid_In(add_kernel52_Valid_Out),
		.Data_Out(bn52_Data_Out),
		.Valid_Out(bn52_Valid_Out)
	);
	Relu_Core rl_kernel52(
		.Data_In(bn52_Data_Out),
		.Valid_In(bn52_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(rl52_Valid_Out)
	);
//////////KERNEL53//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111110101100010011011001111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111101011001011101110010100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111101110001011100101001010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110100011011100111001111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111100100100001101001011000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111101100001010110110010001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111110010100011110000111011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111100111100110100001101110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111101111101010111010101100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111101000101000110000010101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111101010110011101011111000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111110010011001100011101101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111101101110101101101100000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111101110111111011010001010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110011000010010001111011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111101011111000001101100100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110111001011011100010000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111101001111101100010001100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110100000100100001010000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110100100101110100101001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110010001000101101001010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111100101110001001100100110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110011001010011001110011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111110101000100101100010111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111110000111100100001000010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111101111011111001000001001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110011011100101101110101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111110000001010101111010011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111110000110100110100000101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111110011010010111100101010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111110000010110110111000001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110000011111011001000101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b00111100010001010101010000101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b00111101001001010101010011101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111110100010010101111100111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111011100001001110111000101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111110100011000100000100101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111100111111110110010110111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b00111110010101100000101000100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111101110000011011000010110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111111000010000000001010010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111101110000011101011101100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111101101100011001010101001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111101111011101001000000100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111110001110110001001111010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111110100110101111101110000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111110010010011000000100111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111110101000101011011010101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111101001010101100001010010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b00111101000001110101111110111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111110010101011010011001111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111110001100111011101010001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b00111101101010111001011101000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111110110101100111101000001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b10111101011111010111011100010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111101101010010111010101110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111110101101011010001001101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111101000111111101011000111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b10111101101001011011101010010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b00111101101011110011100111010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111110000100001111001010110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b10111010011100011000001011111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111110000110000100000110100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111100010100111110011110111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel53_Valid_Out)
	);
	Adder_64input add_k53(
		.Data1(Data_Out_Kernel53[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel53[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel53[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel53[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel53[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel53[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel53[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel53[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel53[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel53[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel53[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel53[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel53[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel53[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel53[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel53[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel53[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel53[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel53[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel53[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel53[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel53[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel53[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel53[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel53[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel53[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel53[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel53[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel53[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel53[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel53[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel53[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel53[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel53[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel53[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel53[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel53[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel53[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel53[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel53[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel53[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel53[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel53[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel53[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel53[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel53[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel53[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel53[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel53[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel53[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel53[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel53[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel53[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel53[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel53[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel53[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel53[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel53[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel53[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel53[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel53[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel53[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel53[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel53[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel53),
		.Data_Out(add_k53_Data_Out),
		.Valid_Out(add_kernel53_Valid_Out)
	);
	Batch_Norm bn_kernel53(
		.Data_A(32'b00111110011000001100001011011001),
		.Data_B(32'b10111111000001001001100101110000),
		.Data_In(add_k53_Data_Out),
		.Valid_In(add_kernel53_Valid_Out),
		.Data_Out(bn53_Data_Out),
		.Valid_Out(bn53_Valid_Out)
	);
	Relu_Core rl_kernel53(
		.Data_In(bn53_Data_Out),
		.Valid_In(bn53_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(rl53_Valid_Out)
	);
//////////KERNEL54//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110010100110010001001110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111101010000111011011011000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110001011101010000010110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111101111001011010001100110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111110010000101111010100011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110001101100110010001101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111111000111111110010000111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111111010011110110011111111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111110100011101101110100001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110010000110101110111011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111110110101010110001110101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110001100100001111010010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111111001110100010110010100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111110110101001010010110110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111101100101000110001000011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111111001110100110000110010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111100111100010110100111011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111101010100101101000100010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110100100110111001001100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110101110000000110101000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110000000011101010100100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111110110111110110010100101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110111011101001010011000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111110101111100111101101010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111101110100110101110001110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110110101110010001000110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111110111110001101111111101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110111111010110111100111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111111010101101111101011010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110101011010011111111011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111110000111011111110010110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111110010110111100101000000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111110101101011101000011110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b00111101101010110110111001000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111101111111000100111001111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111110100111001100011010000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111101110111011100001101001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111110110101001010010110101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111110101110101001010010101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b00111110000010010010111010000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b10111100101000010001101101101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111100001110000100100010010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b00111110101101010111110001001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b00111110100100010011110101011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111110101011011101001111010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b10111111000000001110010101001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111101110111101110001001101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b00111110101010110110010010101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b00111101001101010000111000011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b00111101100011101010111010101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111110110011000101000000100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b10111001010111001111010101110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111110110101111111110011101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111100011101010011001100010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111110101110010010100101111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b00111111010000001011100100111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b10111110011001110111100110000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111110000001010000111111110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b10111110011010000001110001101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111101010110010001010011001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111110101011001111011011011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111101100000100010101000011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111110101110010100110010110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b10111101010010010100001101110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel54_Valid_Out)
	);
	Adder_64input add_k54(
		.Data1(Data_Out_Kernel54[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel54[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel54[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel54[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel54[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel54[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel54[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel54[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel54[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel54[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel54[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel54[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel54[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel54[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel54[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel54[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel54[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel54[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel54[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel54[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel54[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel54[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel54[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel54[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel54[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel54[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel54[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel54[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel54[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel54[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel54[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel54[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel54[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel54[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel54[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel54[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel54[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel54[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel54[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel54[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel54[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel54[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel54[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel54[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel54[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel54[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel54[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel54[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel54[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel54[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel54[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel54[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel54[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel54[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel54[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel54[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel54[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel54[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel54[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel54[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel54[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel54[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel54[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel54[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel54),
		.Data_Out(add_k54_Data_Out),
		.Valid_Out(add_kernel54_Valid_Out)
	);
	Batch_Norm bn_kernel54(
		.Data_A(32'b00111110010011010011101110100010),
		.Data_B(32'b10111110010101000000100100110110),
		.Data_In(add_k54_Data_Out),
		.Valid_In(add_kernel54_Valid_Out),
		.Data_Out(bn54_Data_Out),
		.Valid_Out(bn54_Valid_Out)
	);
	Relu_Core rl_kernel54(
		.Data_In(bn54_Data_Out),
		.Valid_In(bn54_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(rl54_Valid_Out)
	);
//////////KERNEL55//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111101001111010000011111011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110101010101000001100110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111101000110000110010001101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111111000010010111010100000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111101011110011110100110001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110000001110000001000110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111110100111001101100010001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111110011101000110110111110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110111100101110101111100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111101110101000111000001110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111111001110100010000011100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110100000000000110010110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111110000000100010010000010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111111000010110000111111010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111101111101000001001011111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111110000000111110000101000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111111000011101000111010101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111110101000101010010100011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111110110111001011101110100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110100100011000111011101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110111110110001110010100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111110010001011001000110110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111101001010000010010101110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111111000111101100010101100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111110011111101101001011011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111111001000001000010010010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110010010111001100010100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111110100111001100100001110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111110110111001111000000111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111111000001100001001000101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111100011101001001001000100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111111011111100110000110011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b00111110110010011010011111100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b00111101001001101101100100100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111110010001101110110011010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111101010010011000001010011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111101110000101011101011101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b00111101101111100000011000101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b00111110111000000111100000101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111110101000111001001001001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111111011101000110111010001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111111000001001000110111011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111110000110111101000111000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111110001101001010101000010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111101111000000000000100110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111110000001101010100010111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b10111110001000100011110111011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111110110001000111110010001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b00111100000010100000101100011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b00111110011100110011001011111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b10111011010010100010111111100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111110000001110011110010100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111101110100101000110000000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111110101101101111000101111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b10111110100000110110110011110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111110101000111010000110100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b10111110100100001000110000010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b10111110001011110010010001000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b10111101001000010000010010001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111110101000110110001010010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b10111110010101011010110111100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111110011111010101110101011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111110111000010111101101001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b10111111000000110011010100101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel55_Valid_Out)
	);
	Adder_64input add_k55(
		.Data1(Data_Out_Kernel55[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel55[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel55[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel55[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel55[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel55[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel55[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel55[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel55[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel55[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel55[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel55[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel55[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel55[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel55[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel55[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel55[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel55[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel55[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel55[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel55[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel55[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel55[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel55[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel55[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel55[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel55[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel55[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel55[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel55[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel55[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel55[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel55[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel55[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel55[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel55[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel55[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel55[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel55[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel55[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel55[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel55[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel55[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel55[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel55[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel55[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel55[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel55[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel55[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel55[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel55[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel55[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel55[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel55[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel55[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel55[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel55[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel55[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel55[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel55[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel55[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel55[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel55[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel55[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel55),
		.Data_Out(add_k55_Data_Out),
		.Valid_Out(add_kernel55_Valid_Out)
	);
	Batch_Norm bn_kernel55(
		.Data_A(32'b00111110001000011011100000101001),
		.Data_B(32'b10111110110101000100101000100000),
		.Data_In(add_k55_Data_Out),
		.Valid_In(add_kernel55_Valid_Out),
		.Data_Out(bn55_Data_Out),
		.Valid_Out(bn55_Valid_Out)
	);
	Relu_Core rl_kernel55(
		.Data_In(bn55_Data_Out),
		.Valid_In(bn55_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(rl55_Valid_Out)
	);
//////////KERNEL56//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110100111000110100011110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111110100101001011100010100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110000110111110110100101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111111000101110110000110011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111101011111001001000011010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111100100111011010100010010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111101011101001100101111000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111101000111111000010011101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111110101000100111110111000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110000000000001111111111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111100111001001010100011010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111101000111111001010101100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111100101110111001100110111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111101111001101001011011011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110100111001010001110001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111110011011001111000110101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111111001110010111001001100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111101111100100111110110101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111110101000110001011000000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111110000111001101011110100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110100110000011010111001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111110011011000010100111000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111110101111100110011000000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111110110100110110101100001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111110011011001001111011101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111110111000001011000010000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111110010101001000010011001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111101100010001110100101010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111110011010101010001111110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110000010000101100101010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111110011000110000000001011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111110011101010000001000100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b00111110001011111001101000100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111110100000100010011000000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111111001001011001010010111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111101111100111100010110011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b10111110011011100011100010110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111110001111001011011010100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111110100101000110000001110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b00111010100101100111000000101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b10111110110111110010110110001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b10111101010110011001011010011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111101110111001110100101000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b00111101100111011100101011000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b00111110001111111111101110010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b10111110100000111011100100100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b10111101001100011100101110000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b00111110101100011100010110111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111101100000001111110101001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111100010011001011110001000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111100011110111101011110101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b10111110110110110100000001111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111101010111000101101000101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b00111110010011011100010111110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111110011011011000101110010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111101100011010000100000001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b10111111000100100000011000110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b10111101111100110010000000100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111101101001100010110011111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b00111101110001101101011100100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111101001100111101001011111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b10111110001001101000111001000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b10111100000100001110111100111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111110101010111011100101000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel56_Valid_Out)
	);
	Adder_64input add_k56(
		.Data1(Data_Out_Kernel56[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel56[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel56[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel56[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel56[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel56[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel56[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel56[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel56[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel56[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel56[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel56[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel56[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel56[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel56[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel56[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel56[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel56[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel56[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel56[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel56[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel56[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel56[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel56[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel56[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel56[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel56[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel56[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel56[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel56[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel56[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel56[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel56[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel56[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel56[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel56[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel56[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel56[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel56[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel56[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel56[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel56[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel56[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel56[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel56[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel56[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel56[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel56[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel56[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel56[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel56[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel56[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel56[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel56[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel56[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel56[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel56[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel56[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel56[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel56[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel56[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel56[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel56[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel56[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel56),
		.Data_Out(add_k56_Data_Out),
		.Valid_Out(add_kernel56_Valid_Out)
	);
	Batch_Norm bn_kernel56(
		.Data_A(32'b00111110001101011011111011010011),
		.Data_B(32'b00111111001110000111011010101011),
		.Data_In(add_k56_Data_Out),
		.Valid_In(add_kernel56_Valid_Out),
		.Data_Out(bn56_Data_Out),
		.Valid_Out(bn56_Valid_Out)
	);
	Relu_Core rl_kernel56(
		.Data_In(bn56_Data_Out),
		.Valid_In(bn56_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(rl56_Valid_Out)
	);
//////////KERNEL57//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110100110101011011011100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111111000001010111101011100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110101001010001000111100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111111000010001111101000111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111110011011100100101110100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111110001100100000101001111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111110100101011111000111010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111110010011100111100111101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111101111100100001010000110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111100101001011111100000111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110010011111110100010110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111101101100011011001010110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111101101000011001000101110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111110110000000100100000011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110010011100100011101010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111110110000001101111101001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111110110110010011101000001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110100100101010110011001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110000000000010011000101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111100100011100100000101000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110101001000111110011010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111101101110000011010011011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111111100000100011100001111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111110100010101001100010011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111111000100010111110110011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111110110100001011000101100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110010001011101101011110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111110110001000010010100101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111101101011011011100001110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111101110000110100000100000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111101001010001011011101011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111111000101000110001110000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111100011010011001010111011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111110101101101110110110011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111110110010001111001010001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b10111101110001001011010110000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b10111111010010010010011011001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111110110011110101001110001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111110111000010111101110001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111100101011001111111011010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b10111111001010100100101010100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b10111101111110111011011011100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b00111110011000010111111001100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111110010111111110001011011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b00111110101011111011010111011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b10111110011000000110111011101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b10111110000110101001000010000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b00111101010100110001111101010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b00111110100001010001101101011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111101100101000010110100000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b10111110100101001001111110011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b10111110001011011110111111000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111110010111100101000011110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111101001111000000000110010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111110001101110001111110110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111101001001011010010111001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b10111110101011101111100101110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b10111101011011010010000011010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111101111000111010011000010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b00111110000110001001010011011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b10111110100000100110000110101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b10111101110000110001001111010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b10111110101001001000100101011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111110000001010000000000111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel57_Valid_Out)
	);
	Adder_64input add_k57(
		.Data1(Data_Out_Kernel57[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel57[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel57[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel57[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel57[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel57[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel57[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel57[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel57[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel57[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel57[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel57[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel57[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel57[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel57[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel57[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel57[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel57[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel57[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel57[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel57[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel57[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel57[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel57[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel57[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel57[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel57[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel57[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel57[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel57[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel57[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel57[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel57[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel57[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel57[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel57[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel57[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel57[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel57[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel57[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel57[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel57[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel57[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel57[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel57[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel57[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel57[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel57[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel57[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel57[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel57[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel57[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel57[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel57[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel57[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel57[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel57[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel57[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel57[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel57[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel57[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel57[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel57[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel57[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel57),
		.Data_Out(add_k57_Data_Out),
		.Valid_Out(add_kernel57_Valid_Out)
	);
	Batch_Norm bn_kernel57(
		.Data_A(32'b00111110000100011001100100001011),
		.Data_B(32'b00111111100011100011011111011111),
		.Data_In(add_k57_Data_Out),
		.Valid_In(add_kernel57_Valid_Out),
		.Data_Out(bn57_Data_Out),
		.Valid_Out(bn57_Valid_Out)
	);
	Relu_Core rl_kernel57(
		.Data_In(bn57_Data_Out),
		.Valid_In(bn57_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(rl57_Valid_Out)
	);
//////////KERNEL58//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111110110101001010000011011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110100110011111101001011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111101111100101010101001010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110000011100101100010001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111101110101000100111001110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111101010111110101110101000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111110010111001111101111001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111101001001110011100100100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111101100100110011011011100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111110000011110010000001101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111100011101100101100101001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111101000000101000011100011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111101010010101100001000100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111100011000111011001011101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110011001111101110011100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111110100100011001011111111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110001011100110110101011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110011000001100100110001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110001100011011011010101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111100100001001111100000011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110101010010100000100110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111110011101011100111110001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111101100111101100011011010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111110000111110011010001101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111101011010000111010010001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110101110010111000111111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111111000101110110001101101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110000011100101010101000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111110000110001110111000001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111110100010001100000101000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111110111010101100011100010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110110011000110010001100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b00111101011001111101001000011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b00111110101010000001011111100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111110101111001011010100111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111100100010000010110001010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111101001100010001110000001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111110001011100010100000101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b00111101111101101011001011101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111011111000111110100001000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111111010000010110111001000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111101111001000000001110001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111100101000001111100010010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111110011110000100010010110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111110010100001100110101110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111110110001011110000010011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111110011000111010101010011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111110100000011110000101101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111100011111110011100100100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b00111101100111001011001100100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111101101101000011111001001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111110000101110111111001000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b00111110100100010001111100011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111110101110011010111010011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111101010111111110100011111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111110001111011100001101001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111110100010001000111110000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111110001101111100101101100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b10111110010110010111101011101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b00111100111011010010001011001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111101010101000100011110001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111101111101101001101111101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111111000000000110010101111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b10111110001111101000111101101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel58_Valid_Out)
	);
	Adder_64input add_k58(
		.Data1(Data_Out_Kernel58[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel58[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel58[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel58[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel58[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel58[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel58[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel58[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel58[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel58[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel58[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel58[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel58[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel58[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel58[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel58[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel58[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel58[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel58[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel58[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel58[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel58[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel58[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel58[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel58[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel58[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel58[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel58[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel58[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel58[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel58[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel58[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel58[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel58[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel58[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel58[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel58[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel58[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel58[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel58[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel58[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel58[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel58[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel58[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel58[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel58[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel58[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel58[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel58[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel58[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel58[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel58[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel58[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel58[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel58[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel58[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel58[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel58[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel58[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel58[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel58[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel58[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel58[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel58[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel58),
		.Data_Out(add_k58_Data_Out),
		.Valid_Out(add_kernel58_Valid_Out)
	);
	Batch_Norm bn_kernel58(
		.Data_A(32'b00111110010111100100010010011000),
		.Data_B(32'b10111110101101011011110001110011),
		.Data_In(add_k58_Data_Out),
		.Valid_In(add_kernel58_Valid_Out),
		.Data_Out(bn58_Data_Out),
		.Valid_Out(bn58_Valid_Out)
	);
	Relu_Core rl_kernel58(
		.Data_In(bn58_Data_Out),
		.Valid_In(bn58_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(rl58_Valid_Out)
	);
//////////KERNEL59//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110110111010010000000011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111110110101001110110001101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110011010000001101000011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110110001001010010110001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111101111000100001010111000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111100100010010101000011010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111010000010100010110001100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111101111110001011100110010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111111000010000111010010110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111101111011111010111110100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111101010101010111011000101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111110010010110110000101000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111101100100010001010111010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111101101011010010001011110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110010111000000010010000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111101001001110000010100110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111110110100001010100000100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110100010001100101110000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111101100110110100101101100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111101101000111100110111100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110110000011011011100110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111101010000110110111100011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111110111000001000001111010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111110101010010110100100110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111110101010001011010000011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111110111100111100111111110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111110100001000010000000000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111110111000100111111010010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111110011100110000101001010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110011100010110100010010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111011100100011010110011001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111110101001010010101101110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b00111110010100011101010001100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111100111111111110011011110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111111000010011011000101101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111101111110100111001111100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b10111110110001110100001111011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111110000101000000111100010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111110010000100000100100101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111101111101010100101011100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b10111110110101110110110010001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b10111101101110110101100110000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b00111110000001000000111101110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111110001000100000101011010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b00111110110010010000010110100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b10111110101110101111100110011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111100101110010001011010011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b00111110100111010010000011000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111110000001101000101010010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111101010111100101010100011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b10111101100000101101100000111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b10111110100011111001111100101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111101111001110110010000101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b00111110011010101001111011101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111101100010011000001110000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b00111101101100000100101001001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b10111110111000111111111010101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b10111110010010000000110100101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111101000101010000100010000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111100110010001001101011000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b10111110001010100000001100010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b10111101000011101100000001101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111011111111001011111011100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111101100000001010111011010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel59_Valid_Out)
	);
	Adder_64input add_k59(
		.Data1(Data_Out_Kernel59[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel59[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel59[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel59[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel59[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel59[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel59[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel59[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel59[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel59[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel59[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel59[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel59[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel59[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel59[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel59[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel59[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel59[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel59[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel59[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel59[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel59[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel59[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel59[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel59[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel59[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel59[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel59[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel59[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel59[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel59[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel59[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel59[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel59[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel59[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel59[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel59[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel59[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel59[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel59[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel59[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel59[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel59[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel59[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel59[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel59[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel59[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel59[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel59[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel59[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel59[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel59[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel59[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel59[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel59[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel59[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel59[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel59[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel59[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel59[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel59[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel59[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel59[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel59[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel59),
		.Data_Out(add_k59_Data_Out),
		.Valid_Out(add_kernel59_Valid_Out)
	);
	Batch_Norm bn_kernel59(
		.Data_A(32'b00111110001101111011110110011110),
		.Data_B(32'b00111111010001110000100010110001),
		.Data_In(add_k59_Data_Out),
		.Valid_In(add_kernel59_Valid_Out),
		.Data_Out(bn59_Data_Out),
		.Valid_Out(bn59_Valid_Out)
	);
	Relu_Core rl_kernel59(
		.Data_In(bn59_Data_Out),
		.Valid_In(bn59_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(rl59_Valid_Out)
	);
//////////KERNEL60//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111101110111010010010111111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111110100100011010011111000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111111011001100001101101000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111111010100001110100000011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111101100000100010011101010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111110010000111001010011101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111110110010010010011111101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111100111100101010010011100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111110010011011011000010100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111110010111111101000011110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111111000110100000100000110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111101010011001000110110011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111100110100101000101101001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111111000001110000110101100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110101001000000101001001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111110010101100011111011000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111110101001001010001011110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110110010111011110010101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111110110010100000110011110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111011100011100000010110001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111101001000010111111011000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111101111100100101111101111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111111011111101011000110111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111110111010101101001110000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111110111111110110101101101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111110101010011001101110011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110101011000000001010011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111110011010100000100100100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111110010010110100101010001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111101110100001010001011010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111110101001110001011000010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111110100111111001001011111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111110011111011100000011011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111100110001001011110100101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111101101110010110110001000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b10111101110110001100010110100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b10111111010011101101100110111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111110011101010101110010110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111111001011001001000000010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111101100010110010001011000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b10111111001001000100010001110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111101101110110011110001000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b00111110101001001111000101100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111110101110100111101011010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111101101110110111111111110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b10111110000110100011101000101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111110001010100101111100011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111110001110111100010000101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b00111101111011000101110011011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b00111110010010001110001111001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b10111110010011000011100101111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b10111110011010110011011011001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111110010010111111000011010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b00111101101100100001010110001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111101010010101010001100111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b00111110100101011001110100110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b10111110110110110100100011011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b10111110010101110110111010001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b10111100111111010100100000011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111110100100010110011100010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b10111110001010101010010101010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111101000101011101000000110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b10111111001100001001100010001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111110010111011010110011001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel60_Valid_Out)
	);
	Adder_64input add_k60(
		.Data1(Data_Out_Kernel60[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel60[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel60[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel60[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel60[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel60[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel60[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel60[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel60[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel60[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel60[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel60[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel60[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel60[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel60[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel60[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel60[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel60[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel60[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel60[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel60[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel60[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel60[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel60[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel60[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel60[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel60[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel60[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel60[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel60[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel60[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel60[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel60[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel60[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel60[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel60[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel60[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel60[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel60[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel60[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel60[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel60[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel60[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel60[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel60[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel60[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel60[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel60[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel60[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel60[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel60[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel60[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel60[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel60[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel60[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel60[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel60[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel60[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel60[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel60[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel60[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel60[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel60[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel60[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel60),
		.Data_Out(add_k60_Data_Out),
		.Valid_Out(add_kernel60_Valid_Out)
	);
	Batch_Norm bn_kernel60(
		.Data_A(32'b00111110000100010000011000100100),
		.Data_B(32'b00111111101010000000110101100000),
		.Data_In(add_k60_Data_Out),
		.Valid_In(add_kernel60_Valid_Out),
		.Data_Out(bn60_Data_Out),
		.Valid_Out(bn60_Valid_Out)
	);
	Relu_Core rl_kernel60(
		.Data_In(bn60_Data_Out),
		.Valid_In(bn60_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(rl60_Valid_Out)
	);
//////////KERNEL61//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110111111111110101000111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111101110011010001111011010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110000110110100100110111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110000011110110111110100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111110001100100111010101011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111110011101111111100101101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111110111001101011011110001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111101000101101111000000111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111100001111010101000010110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111100001010111001100101111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111110110011010000110011011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111111000101100100111100100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111100110110001001000001100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111110011011101111100011110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111101111001011110010100011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111110000101000010100001100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111110110101000110011011100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111100001010111001101011100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111110100010000111110101011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111101101000001110010011001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111101111010010011110011100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111110110110101010011111110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111101101110110011110000011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111111000100000010001110100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111110011001110000000100100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111110111100011101000000100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111110000110011000101001010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110101101011010101110011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111110101001001000110000010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110101011111001100010110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111110101001001101110001011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111110110011011100001001010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111110110011001000101001110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b00111110101001001111101100111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111101100111001010001001001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b10111110001111000100101001000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b10111101101001101110011111010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111111000001101111011001100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111111011010100101110111011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b00111110001000111000100000001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b10111111100100110110011101111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b10111111000000000000111000100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b00111101000101100011010111100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111110100111011100100010101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111100100100000000000100110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b10111111000001010010011110110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111110001110011001111111111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b00111110010010110100111101001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111101100101101110101101010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b00111110100101011110010111001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b10111110100110010101001111000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b10111110010001101000011100110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b00111110110000000101010110111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b00111110010001100001101000111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b10111110100110101101011110010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111110010001101000111111101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b10111110101001010111111010000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b10111110100110110010001100010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b10111101100000111011001110001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111101110101011111111011000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b10111110110000111100100010001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b10111110011111100001100000000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b10111111001001001111001101110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111111000101010110110010000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel61_Valid_Out)
	);
	Adder_64input add_k61(
		.Data1(Data_Out_Kernel61[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel61[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel61[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel61[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel61[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel61[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel61[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel61[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel61[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel61[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel61[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel61[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel61[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel61[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel61[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel61[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel61[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel61[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel61[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel61[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel61[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel61[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel61[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel61[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel61[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel61[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel61[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel61[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel61[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel61[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel61[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel61[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel61[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel61[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel61[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel61[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel61[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel61[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel61[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel61[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel61[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel61[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel61[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel61[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel61[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel61[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel61[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel61[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel61[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel61[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel61[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel61[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel61[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel61[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel61[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel61[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel61[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel61[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel61[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel61[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel61[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel61[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel61[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel61[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel61),
		.Data_Out(add_k61_Data_Out),
		.Valid_Out(add_kernel61_Valid_Out)
	);
	Batch_Norm bn_kernel61(
		.Data_A(32'b00111110000110101101011100011100),
		.Data_B(32'b00111111110110001110000011001001),
		.Data_In(add_k61_Data_Out),
		.Valid_In(add_kernel61_Valid_Out),
		.Data_Out(bn61_Data_Out),
		.Valid_Out(bn61_Valid_Out)
	);
	Relu_Core rl_kernel61(
		.Data_In(bn61_Data_Out),
		.Valid_In(bn61_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(rl61_Valid_Out)
	);
//////////KERNEL62//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110111000101001100010010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111110010110000010111100101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111101100101010010111010100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110001001000011010011100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111110001011111111111000111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111101001111110010000001101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111100111001000001111110111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111101100100110000111000001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111111000000101111000010011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110010010110011010000111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110010100101011111011010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111100110110011010101011011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111101111010010000011001001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111110100101110011001011100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110011011100001001011100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111101101100000000100101010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111110100110010001111001111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111101001111110000010110110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111101010101001110011110000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111101011110000000101011000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110110011011101010100110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111101110011110000101100110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111110101010100110111011101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111110000010100000001000011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111110101001010000000101001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111110100110100111000001011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111110110011110111100011011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111111000001111000101101100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111100111110110000000101110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110001101110000010000101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111110000101000000001001010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111110000101001110110100010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b00111110110000001100100001100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111110110100010010110010010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111111001110001011000101110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111101111101111000001111011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b10111110100010011001110111100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111101110100001101100000000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111110100001011010100000001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111101001011011000000010110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b10111110100011101011111000110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b10111101101100011100111010000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b00111101100001011101001101000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111110001100101001101011101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b00111110110011110011111100110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b10111110001010011101000010101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b10111110011010101101101101000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b00111110110101001110001011001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b00111100001010111110001000100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b00111101111001110111001010011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111110011111010100010100010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b10111110011011000111101100010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111110010101000111101000001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b00111110101001100101011111001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b10111101011110000110101101100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b00111101011000001001101010110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b10111110111100011000000111010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b10111110101111101010110111101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111110111010000001110110001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111101111000010110101100010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b10111011101101110001100100010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111101100001100111110101011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111101001101000101000000100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111110000000011101001001111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel62_Valid_Out)
	);
	Adder_64input add_k62(
		.Data1(Data_Out_Kernel62[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel62[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel62[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel62[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel62[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel62[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel62[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel62[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel62[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel62[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel62[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel62[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel62[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel62[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel62[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel62[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel62[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel62[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel62[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel62[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel62[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel62[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel62[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel62[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel62[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel62[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel62[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel62[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel62[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel62[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel62[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel62[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel62[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel62[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel62[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel62[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel62[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel62[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel62[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel62[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel62[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel62[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel62[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel62[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel62[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel62[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel62[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel62[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel62[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel62[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel62[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel62[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel62[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel62[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel62[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel62[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel62[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel62[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel62[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel62[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel62[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel62[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel62[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel62[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel62),
		.Data_Out(add_k62_Data_Out),
		.Valid_Out(add_kernel62_Valid_Out)
	);
	Batch_Norm bn_kernel62(
		.Data_A(32'b00111110010000101110100011101010),
		.Data_B(32'b00111101111010110101001101110000),
		.Data_In(add_k62_Data_Out),
		.Valid_In(add_kernel62_Valid_Out),
		.Data_Out(bn62_Data_Out),
		.Valid_Out(bn62_Valid_Out)
	);
	Relu_Core rl_kernel62(
		.Data_In(bn62_Data_Out),
		.Valid_In(bn62_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(rl62_Valid_Out)
	);
//////////KERNEL63//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111101110010001000101100110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111110101100011100010110000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110110110101010110001010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110110011101001101100001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111101101000110100001011010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111110110000000100100101011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111111001011011010111000100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111110100001110011001011111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111011101101111101100010100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110000011100111101000101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111101101101101110011001111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111101110100110010010010110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111100110101011101001100100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111111001101101011110000010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111101100011011000111101100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111110001110100011101010010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111101110101010100000001100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110101110110101000000000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110000101001111011010111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111101001001001111011010001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110100000001001111101100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111110100011111100111010101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111111010000010100111000110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111101001010001100111110111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111110110000110111000011100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111110110101010100100110010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111101101101111110100101011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111110100011001000000111100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111101010111110001011001000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110101001010101110110111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111101010100010011101111000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111111011100010001111001101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111110110110111101011011001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111110100010001011000100010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111111000010101110101001101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b10111011110111011000111110010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b10111111010111010011101000010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111110111110000100000101111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111111001001110110100000100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b00111110100001001000001111101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b10111110010101111000100001101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b10111110010101110111001000000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b00111110001011100010010100000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111110100001111110101111000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b00111110110001010111010011011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b10111100110010001110100110010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111110100000001011010110110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b00111011101010001110111010001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b00111110110001000000101010000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111101100101000011111101000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b10111110011011100010100110110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b10111110011011001110111000110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111110110111000000100010100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111110010111011000110011101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111110100110101101111001001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b00111110011011011001000001001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b10111110101100100101001111100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111110000111010111011010100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b10111110001100100110001011010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b00111110100011111110000001001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b10111110000100101001000001100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b10111110001101011100001001001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b10111110111010011101100100001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111111000010010111100000011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel63_Valid_Out)
	);
	Adder_64input add_k63(
		.Data1(Data_Out_Kernel63[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel63[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel63[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel63[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel63[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel63[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel63[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel63[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel63[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel63[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel63[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel63[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel63[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel63[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel63[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel63[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel63[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel63[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel63[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel63[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel63[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel63[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel63[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel63[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel63[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel63[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel63[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel63[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel63[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel63[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel63[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel63[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel63[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel63[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel63[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel63[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel63[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel63[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel63[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel63[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel63[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel63[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel63[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel63[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel63[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel63[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel63[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel63[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel63[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel63[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel63[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel63[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel63[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel63[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel63[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel63[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel63[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel63[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel63[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel63[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel63[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel63[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel63[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel63[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel63),
		.Data_Out(add_k63_Data_Out),
		.Valid_Out(add_kernel63_Valid_Out)
	);
	Batch_Norm bn_kernel63(
		.Data_A(32'b00111110001000000001100100010001),
		.Data_B(32'b00111111010110100110001111110101),
		.Data_In(add_k63_Data_Out),
		.Valid_In(add_kernel63_Valid_Out),
		.Data_Out(bn63_Data_Out),
		.Valid_Out(bn63_Valid_Out)
	);
	Relu_Core rl_kernel63(
		.Data_In(bn63_Data_Out),
		.Valid_In(bn63_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(rl63_Valid_Out)
	);
//////////KERNEL64//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110001011011111000111000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111101100011000011100010100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110100100100001010000111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111101001000010001110011011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111101000011110110011100101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110011010011110000101000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111110111100010110011000101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111011110000110100000011111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111110100011001011111000100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111110010111001011101010110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111101111111100101111001001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111110101111011101010101011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111101010001110100100110110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111110110001001110010000011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110011100111110001010011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111101011110000000011010010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110100010101100111010010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111100010001001011110011001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111111000111111111110010110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111110111100111010110000101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111111000110011000001001000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111100110111110100011011001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111100101100111011101011110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111110000001000100101000111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111111000011100111010000111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110100010011111010110101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111111001100100001000111101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111101100011000011111100011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111101010010010000101100100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111111011111110100000101001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111110100001100010001011110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110110110101000000001101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111111000101111111110000111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b00111110110010111110100111011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111110011100011101001001100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b10111110001101001111011111011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111111000011010110100000111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b00111111001101101000101110100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b00111110110010110100111000010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111110101111100000111010111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b10111101001011110111111001101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111111000011001000001010110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b00111101100111100111011101010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b00111110011001010110100110011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111111001010100110110101000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b10111110010010001100110001011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b10111101101001001100100110000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111110100110000100001000000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111111000000101010000001001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b00111110111110001110110110000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111110001010111011110101001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b10111010001101000101110110011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b00111110100010000011110111010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111101101010010110100010010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b10111110101000110101000001000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b00111110011000001100101111101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111101010011010100100111000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b10111110000011101010010010111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111110010010101101110111000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111111010000001001010100000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b10111100100010110100011001000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b10111110000100101000111000010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111110001011111000111100110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111110011000101111111111110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel64_Valid_Out)
	);
	Adder_64input add_k64(
		.Data1(Data_Out_Kernel64[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel64[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel64[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel64[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel64[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel64[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel64[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel64[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel64[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel64[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel64[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel64[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel64[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel64[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel64[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel64[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel64[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel64[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel64[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel64[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel64[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel64[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel64[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel64[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel64[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel64[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel64[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel64[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel64[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel64[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel64[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel64[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel64[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel64[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel64[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel64[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel64[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel64[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel64[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel64[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel64[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel64[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel64[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel64[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel64[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel64[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel64[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel64[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel64[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel64[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel64[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel64[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel64[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel64[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel64[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel64[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel64[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel64[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel64[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel64[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel64[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel64[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel64[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel64[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel64),
		.Data_Out(add_k64_Data_Out),
		.Valid_Out(add_kernel64_Valid_Out)
	);
	Batch_Norm bn_kernel64(
		.Data_A(32'b00111110001101101011000110101100),
		.Data_B(32'b00111111000010011100010000110011),
		.Data_In(add_k64_Data_Out),
		.Valid_In(add_kernel64_Valid_Out),
		.Data_Out(bn64_Data_Out),
		.Valid_Out(bn64_Valid_Out)
	);
	Relu_Core rl_kernel64(
		.Data_In(bn64_Data_Out),
		.Valid_In(bn64_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(rl64_Valid_Out)
	);
//////////KERNEL65//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel65 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110101101010000011011011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel65[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel65_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel65 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111111000111000100010011100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel65[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel65_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel65 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110100011100110100010101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel65[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel65_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel65 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110110100110001111111110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel65[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel65_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel65 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111101111101110010111100011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel65[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel65_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel65 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111011101100001011001001000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel65[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel65_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel65 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111110010101000001101100001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel65[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel65_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel65 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111101001011001000011010010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel65[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel65_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel65 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111110010111110011000001000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel65[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel65_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel65 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110100010001101001101001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel65[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel65_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel65 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110000100111111110001001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel65[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel65_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel65 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110001001000100011000101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel65[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel65_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel65 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111101111000000111111101010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel65[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel65_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel65 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111101100111110110001011010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel65[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel65_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel65 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110101111001011011000110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel65[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel65_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel65 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111100111111110111000100101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel65[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel65_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel65 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111110111011100000001110000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel65[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel65_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel65 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111101000011100101001111110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel65[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel65_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel65 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111101100100011000111100100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel65[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel65_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel65 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111101100100000111011000000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel65[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel65_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel65 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110010111000001001011010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel65[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel65_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel65 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111101100110111010100011111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel65[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel65_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel65 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111110111101111111110011101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel65[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel65_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel65 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111110100001101111000010010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel65[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel65_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel65 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111100110110110111110011110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel65[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel65_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel65 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111110100101000011100001001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel65[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel65_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel65 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111110101101000001101000101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel65[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel65_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel65 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111110100011000101001010010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel65[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel65_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel65 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111110010000011001100001001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel65[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel65_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel65 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110001101001010011001001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel65[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel65_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel65 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111101011111110001010110101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel65[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel65_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel65 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111110111011111010011011010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel65[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel65_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel65 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b00111101001110100010111000111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel65[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel65_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel65 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111110101100101000101111010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel65[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel65_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel65 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111110110000111110111010111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel65[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel65_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel65 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111110000110100100000101111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel65[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel65_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel65 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b10111110100000111101010111011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel65[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel65_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel65 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111101011111101010000011101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel65[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel65_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel65 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111110100000110101001110000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel65[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel65_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel65 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b00111100111100100110010010010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel65[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel65_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel65 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b10111111001111111100100000000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel65[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel65_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel65 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111100100101000100000000100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel65[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel65_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel65 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b00111101010000111000110101101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel65[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel65_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel65 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b00111101000011010110100000011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel65[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel65_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel65 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b00111110010101011111101010110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel65[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel65_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel65 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b10111110101010110111000111000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel65[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel65_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel65 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b10111110000000101110101101000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel65[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel65_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel65 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b00111110100110011000001101000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel65[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel65_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel65 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b00111101000101100101001110111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel65[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel65_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel65 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111101011001101001110001000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel65[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel65_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel65 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111101011100010001011000001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel65[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel65_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel65 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b10111110101010011011101101011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel65[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel65_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel65 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111110100101100100100101010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel65[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel65_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel65 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111101000011100111101111011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel65[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel65_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel65 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111101011111101101111000111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel65[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel65_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel65 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111110000101110101110011001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel65[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel65_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel65 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b10111110011111101110010101110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel65[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel65_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel65 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b10111110111001010101110111101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel65[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel65_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel65 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111110001010111110110011100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel65[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel65_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel65 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111101110011001010001001011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel65[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel65_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel65 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b10111110001110010101010110000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel65[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel65_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel65 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111101010001001011011111001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel65[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel65_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel65 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b10111110000100010100000111110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel65[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel65_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel65 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111110010111010001101000000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel65[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel65_Valid_Out)
	);
	Adder_64input add_k65(
		.Data1(Data_Out_Kernel65[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel65[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel65[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel65[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel65[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel65[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel65[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel65[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel65[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel65[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel65[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel65[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel65[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel65[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel65[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel65[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel65[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel65[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel65[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel65[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel65[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel65[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel65[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel65[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel65[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel65[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel65[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel65[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel65[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel65[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel65[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel65[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel65[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel65[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel65[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel65[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel65[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel65[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel65[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel65[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel65[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel65[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel65[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel65[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel65[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel65[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel65[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel65[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel65[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel65[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel65[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel65[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel65[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel65[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel65[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel65[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel65[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel65[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel65[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel65[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel65[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel65[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel65[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel65[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel65),
		.Data_Out(add_k65_Data_Out),
		.Valid_Out(add_kernel65_Valid_Out)
	);
	Batch_Norm bn_kernel65(
		.Data_A(32'b00111110001101110010110011000101),
		.Data_B(32'b00111111010010110010110010100010),
		.Data_In(add_k65_Data_Out),
		.Valid_In(add_kernel65_Valid_Out),
		.Data_Out(bn65_Data_Out),
		.Valid_Out(bn65_Valid_Out)
	);
	Relu_Core rl_kernel65(
		.Data_In(bn65_Data_Out),
		.Valid_In(bn65_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*65-1:DATA_WIDHT*64]),
		.Valid_Out(rl65_Valid_Out)
	);
//////////KERNEL66//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel66 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110001100010001100100000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel66[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel66_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel66 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111110110111010000100100111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel66[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel66_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel66 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110011110000100101000101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel66[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel66_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel66 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110101101110100111011010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel66[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel66_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel66 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111110001001111111100011100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel66[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel66_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel66 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111101011101000001100110110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel66[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel66_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel66 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111110110001100100011001100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel66[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel66_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel66 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111010110011100100001001101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel66[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel66_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel66 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111110100110010010101100110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel66[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel66_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel66 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111101100000101101100000110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel66[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel66_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel66 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111101111100111110010100100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel66[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel66_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel66 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110010001000111001111111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel66[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel66_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel66 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111100110000000101000010101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel66[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel66_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel66 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111101101111001100110111010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel66[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel66_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel66 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110101010011001001000011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel66[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel66_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel66 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111101101110110111000110000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel66[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel66_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel66 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111111000111001101101111100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel66[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel66_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel66 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111110010001111101000111010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel66[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel66_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel66 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111100101110110010111001001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel66[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel66_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel66 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111100110100100100011001001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel66[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel66_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel66 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110100001001110101010111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel66[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel66_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel66 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111100001101000101111000100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel66[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel66_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel66 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111110100100111111111000011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel66[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel66_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel66 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111110100101010001010111010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel66[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel66_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel66 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111100010111010011001011011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel66[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel66_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel66 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111101111011100001111001010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel66[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel66_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel66 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111110101000111010010010100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel66[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel66_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel66 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111110001011111111100101011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel66[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel66_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel66 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111101001111100010101011000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel66[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel66_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel66 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110110110110100000011010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel66[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel66_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel66 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111110010110011010001000111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel66[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel66_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel66 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111110101111000000100000011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel66[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel66_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel66 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b00111100000011000011001111011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel66[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel66_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel66 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111110100101000000010100111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel66[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel66_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel66 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111110001110001001001101000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel66[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel66_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel66 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111101100011101001001111011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel66[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel66_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel66 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b10111110101111000101110101111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel66[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel66_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel66 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b00111101111001011110111001011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel66[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel66_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel66 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111110101111101110011010110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel66[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel66_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel66 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b00111110011101001110000100110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel66[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel66_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel66 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b10111111011100100111111111000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel66[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel66_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel66 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111101001101100010001110001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel66[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel66_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel66 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b00111110010010110110011111101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel66[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel66_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel66 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b00111110010010111110010111011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel66[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel66_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel66 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b00111110110100000011000001010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel66[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel66_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel66 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b10111101111111000111110101101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel66[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel66_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel66 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b10111110011100100101011010101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel66[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel66_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel66 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b00111110000111001010011111001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel66[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel66_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel66 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b00111101001101111111110110110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel66[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel66_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel66 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111110010001110110111100001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel66[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel66_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel66 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111010110111101111001110100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel66[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel66_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel66 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b10111110011101110110101111000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel66[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel66_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel66 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111110011000111001011100010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel66[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel66_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel66 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b00111101000001001000100110000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel66[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel66_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel66 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111010100101101001101001111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel66[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel66_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel66 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111110000010101110100110110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel66[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel66_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel66 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b10111110010110111010111100000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel66[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel66_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel66 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b10111110101111011111001111000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel66[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel66_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel66 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111101111000001110011101110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel66[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel66_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel66 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111110001001111001101111110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel66[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel66_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel66 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b10111101101010011001100001001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel66[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel66_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel66 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111101100001011100111111010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel66[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel66_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel66 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b10111110101110000110001000011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel66[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel66_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel66 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111110001111111101111001001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel66[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel66_Valid_Out)
	);
	Adder_64input add_k66(
		.Data1(Data_Out_Kernel66[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel66[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel66[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel66[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel66[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel66[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel66[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel66[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel66[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel66[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel66[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel66[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel66[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel66[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel66[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel66[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel66[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel66[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel66[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel66[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel66[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel66[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel66[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel66[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel66[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel66[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel66[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel66[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel66[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel66[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel66[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel66[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel66[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel66[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel66[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel66[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel66[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel66[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel66[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel66[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel66[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel66[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel66[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel66[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel66[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel66[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel66[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel66[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel66[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel66[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel66[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel66[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel66[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel66[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel66[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel66[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel66[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel66[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel66[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel66[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel66[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel66[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel66[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel66[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel66),
		.Data_Out(add_k66_Data_Out),
		.Valid_Out(add_kernel66_Valid_Out)
	);
	Batch_Norm bn_kernel66(
		.Data_A(32'b00111110001010110001101001010001),
		.Data_B(32'b00111110100110001101011000010111),
		.Data_In(add_k66_Data_Out),
		.Valid_In(add_kernel66_Valid_Out),
		.Data_Out(bn66_Data_Out),
		.Valid_Out(bn66_Valid_Out)
	);
	Relu_Core rl_kernel66(
		.Data_In(bn66_Data_Out),
		.Valid_In(bn66_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*66-1:DATA_WIDHT*65]),
		.Valid_Out(rl66_Valid_Out)
	);
//////////KERNEL67//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel67 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111111000000111011001010011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel67[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel67_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel67 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111101010001110000000000101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel67[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel67_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel67 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110000000010011011001110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel67[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel67_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel67 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110000010100100101100010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel67[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel67_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel67 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111101111001010100110111000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel67[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel67_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel67 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111101011001010100011110000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel67[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel67_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel67 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111110010010101100001011100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel67[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel67_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel67 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111101010101011011111101100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel67[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel67_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel67 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110010110111011010011011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel67[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel67_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel67 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111101101110100100111111011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel67[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel67_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel67 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111101110001101101000101110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel67[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel67_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel67 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111101111111100010100101011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel67[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel67_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel67 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110001100000101101000101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel67[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel67_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel67 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111101110001100001110010010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel67[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel67_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel67 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110010011110111010111010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel67[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel67_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel67 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111101100011101101010010000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel67[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel67_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel67 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110100011101101110001010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel67[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel67_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel67 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111101011111101000110011110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel67[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel67_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel67 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110001010110010011000011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel67[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel67_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel67 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110011110111111100010000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel67[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel67_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel67 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110100010101000000101010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel67[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel67_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel67 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111011001101111101011101011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel67[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel67_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel67 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110100110110001010110100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel67[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel67_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel67 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111101111011111110000000110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel67[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel67_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel67 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111110011000110001100011110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel67[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel67_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel67 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110100000010011110110101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel67[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel67_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel67 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110100110000110110100011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel67[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel67_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel67 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110010000011100100100101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel67[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel67_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel67 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111101110110010111100010101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel67[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel67_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel67 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111110001111011101000100000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel67[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel67_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel67 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111110100000011110111000110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel67[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel67_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel67 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111101100011100011110100100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel67[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel67_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel67 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111110010011111110010000100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel67[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel67_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel67 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b00111110100011001001111000110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel67[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel67_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel67 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111110110101011000110011100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel67[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel67_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel67 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b10111101111100001100110001110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel67[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel67_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel67 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111110110011011111000001000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel67[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel67_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel67 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111101101001100110100100000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel67[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel67_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel67 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111100101101100101001101010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel67[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel67_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel67 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111101100001111000001011110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel67[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel67_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel67 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111110111011100101111011001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel67[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel67_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel67 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111110000010001110001000000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel67[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel67_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel67 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111101101011000001011010001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel67[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel67_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel67 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111101101101111011101010000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel67[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel67_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel67 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111110001011111000111110001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel67[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel67_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel67 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111110101011001000000110010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel67[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel67_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel67 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111110110000001100111110010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel67[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel67_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel67 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111110101001001110001000011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel67[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel67_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel67 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b00111101100001111111011111101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel67[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel67_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel67 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111100010000010011101000001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel67[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel67_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel67 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111101111110010110110010011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel67[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel67_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel67 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111110010110010100000001101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel67[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel67_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel67 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b00111101010111111110110101000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel67[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel67_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel67 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111110111101000111000100001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel67[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel67_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel67 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111101111011000111001011001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel67[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel67_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel67 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111110010100100110001110111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel67[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel67_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel67 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111110110011101101101011110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel67[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel67_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel67 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111110000010110101100100001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel67[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel67_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel67 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b10111110000111001011100001011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel67[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel67_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel67 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b00111110000000000111111000001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel67[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel67_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel67 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111101101011101110101100010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel67[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel67_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel67 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111010101011110001000110010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel67[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel67_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel67 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111100011001001100111011111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel67[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel67_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel67 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111100000001000011011111101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel67[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel67_Valid_Out)
	);
	Adder_64input add_k67(
		.Data1(Data_Out_Kernel67[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel67[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel67[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel67[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel67[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel67[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel67[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel67[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel67[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel67[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel67[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel67[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel67[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel67[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel67[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel67[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel67[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel67[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel67[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel67[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel67[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel67[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel67[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel67[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel67[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel67[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel67[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel67[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel67[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel67[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel67[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel67[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel67[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel67[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel67[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel67[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel67[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel67[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel67[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel67[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel67[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel67[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel67[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel67[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel67[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel67[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel67[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel67[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel67[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel67[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel67[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel67[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel67[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel67[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel67[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel67[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel67[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel67[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel67[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel67[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel67[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel67[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel67[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel67[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel67),
		.Data_Out(add_k67_Data_Out),
		.Valid_Out(add_kernel67_Valid_Out)
	);
	Batch_Norm bn_kernel67(
		.Data_A(32'b00111110011000101100101100101100),
		.Data_B(32'b10111110110111010001100010100000),
		.Data_In(add_k67_Data_Out),
		.Valid_In(add_kernel67_Valid_Out),
		.Data_Out(bn67_Data_Out),
		.Valid_Out(bn67_Valid_Out)
	);
	Relu_Core rl_kernel67(
		.Data_In(bn67_Data_Out),
		.Valid_In(bn67_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*67-1:DATA_WIDHT*66]),
		.Valid_Out(rl67_Valid_Out)
	);
//////////KERNEL68//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel68 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111101111100100000101101100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel68[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel68_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel68 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110101011111010000101000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel68[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel68_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel68 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110000100011110111001011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel68[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel68_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel68 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111101100110110011010111111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel68[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel68_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel68 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111110101011011000011010101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel68[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel68_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel68 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111101101100001110001101111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel68[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel68_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel68 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111110101010111001000001101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel68[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel68_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel68 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111011101110001001001000110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel68[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel68_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel68 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111111001110110110111010100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel68[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel68_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel68 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111110000001100010110100010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel68[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel68_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel68 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111111001011001111111110111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel68[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel68_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel68 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111100110111111000011110111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel68[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel68_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel68 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110000010111101111101101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel68[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel68_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel68 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111110001000001110101011111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel68[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel68_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel68 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111101100110010001011100100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel68[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel68_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel68 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111101011011000111010000001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel68[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel68_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel68 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111111000101101110110010001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel68[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel68_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel68 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111101111010001100110001001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel68[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel68_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel68 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111111000111110001111000001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel68[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel68_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel68 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110100100100011000010001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel68[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel68_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel68 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110101001011011101110000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel68[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel68_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel68 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111110001100100000011110011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel68[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel68_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel68 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111011111010001011001000111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel68[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel68_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel68 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111111001000101110111011011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel68[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel68_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel68 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111110001101001001100010000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel68[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel68_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel68 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111100011001100100000110000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel68[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel68_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel68 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111111000111001001011110110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel68[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel68_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel68 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110100100010100010001100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel68[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel68_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel68 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111111000110010111011000001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel68[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel68_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel68 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110101010000011100001101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel68[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel68_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel68 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111110100011010010001111001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel68[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel68_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel68 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110100110111101100100101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel68[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel68_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel68 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111111000001110011110100111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel68[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel68_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel68 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b00111110110101010000100011000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel68[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel68_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel68 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111110110111111010111101100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel68[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel68_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel68 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111010011010010101000011111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel68[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel68_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel68 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111110111011101111011001111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel68[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel68_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel68 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111110011010110001111101110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel68[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel68_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel68 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b00111110010010101111101101111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel68[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel68_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel68 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111001111111010101001010110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel68[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel68_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel68 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111111001000000010111100000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel68[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel68_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel68 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b10111101110111010000010001010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel68[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel68_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel68 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111101101010010010100100010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel68[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel68_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel68 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111101101110010110110000110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel68[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel68_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel68 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111110100010101011100111011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel68[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel68_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel68 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111111000010000011110100010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel68[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel68_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel68 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111110100001101100110100110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel68[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel68_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel68 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111110111110100010001101001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel68[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel68_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel68 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111110011110101111011001010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel68[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel68_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel68 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b00111101100010011000000110001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel68[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel68_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel68 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b10111100110111000010011000111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel68[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel68_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel68 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111110111011111101001110111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel68[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel68_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel68 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b00111101011010001101011110001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel68[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel68_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel68 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111110110110100010010100011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel68[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel68_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel68 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b10111101101100101101001100101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel68[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel68_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel68 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111111001000000111011100010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel68[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel68_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel68 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b10111101111101001000101010010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel68[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel68_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel68 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b10111101010111111000111000110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel68[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel68_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel68 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b10111110010001100100100010101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel68[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel68_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel68 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b00111110011011010101010000100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel68[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel68_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel68 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b10111101101100001111101011011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel68[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel68_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel68 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111110011100000001111100010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel68[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel68_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel68 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111100111111011100110110100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel68[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel68_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel68 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111110000100011100010101000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel68[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel68_Valid_Out)
	);
	Adder_64input add_k68(
		.Data1(Data_Out_Kernel68[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel68[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel68[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel68[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel68[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel68[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel68[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel68[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel68[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel68[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel68[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel68[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel68[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel68[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel68[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel68[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel68[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel68[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel68[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel68[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel68[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel68[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel68[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel68[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel68[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel68[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel68[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel68[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel68[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel68[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel68[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel68[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel68[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel68[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel68[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel68[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel68[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel68[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel68[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel68[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel68[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel68[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel68[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel68[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel68[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel68[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel68[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel68[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel68[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel68[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel68[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel68[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel68[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel68[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel68[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel68[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel68[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel68[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel68[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel68[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel68[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel68[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel68[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel68[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel68),
		.Data_Out(add_k68_Data_Out),
		.Valid_Out(add_kernel68_Valid_Out)
	);
	Batch_Norm bn_kernel68(
		.Data_A(32'b00111110000101101111111011010100),
		.Data_B(32'b10111100000100001010100010101110),
		.Data_In(add_k68_Data_Out),
		.Valid_In(add_kernel68_Valid_Out),
		.Data_Out(bn68_Data_Out),
		.Valid_Out(bn68_Valid_Out)
	);
	Relu_Core rl_kernel68(
		.Data_In(bn68_Data_Out),
		.Valid_In(bn68_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*68-1:DATA_WIDHT*67]),
		.Valid_Out(rl68_Valid_Out)
	);
//////////KERNEL69//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel69 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111110101101101001101111111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel69[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel69_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel69 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110000001000111011101000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel69[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel69_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel69 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110101011100111011001100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel69[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel69_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel69 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110001100010101001010000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel69[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel69_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel69 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111101011101111110000001110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel69[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel69_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel69 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110001001010000101000011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel69[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel69_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel69 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111101000011010011010111000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel69[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel69_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel69 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111110011001101001111011000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel69[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel69_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel69 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111110010000101000001011110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel69[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel69_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel69 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111110011001011101000110110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel69[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel69_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel69 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110000011101010010000111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel69[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel69_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel69 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110000000100101100110001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel69[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel69_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel69 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111101011111001111001111111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel69[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel69_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel69 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111110100011100111000000101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel69[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel69_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel69 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111101110100100011111001100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel69[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel69_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel69 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111101101100110110100011110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel69[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel69_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel69 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111110000011001101011100111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel69[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel69_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel69 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110011100111001101011101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel69[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel69_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel69 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111101000010101100011101000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel69[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel69_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel69 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111101010000011100001111010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel69[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel69_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel69 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110110000010011011110010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel69[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel69_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel69 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111101111010110101111110001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel69[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel69_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel69 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110101010010110000000010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel69[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel69_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel69 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111101111000010001110101011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel69[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel69_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel69 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111101100111000111100111110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel69[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel69_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel69 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110100001101000011100101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel69[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel69_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel69 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111111000100101000001001011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel69[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel69_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel69 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110011111010100011001111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel69[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel69_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel69 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111110001111101010111111010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel69[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel69_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel69 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111110110001001100001111010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel69[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel69_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel69 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111110101110101110001001100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel69[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel69_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel69 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110101110001100010010010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel69[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel69_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel69 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111101110010111101111100011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel69[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel69_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel69 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b00111110100000001011111010101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel69[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel69_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel69 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111111000010000100100100111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel69[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel69_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel69 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b10111110100011010100001110011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel69[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel69_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel69 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111101110110000010000011101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel69[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel69_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel69 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111110001001101111111000101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel69[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel69_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel69 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b00111110000000100110100111100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel69[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel69_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel69 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b00111101000011101110011100100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel69[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel69_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel69 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111111000101000101011100010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel69[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel69_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel69 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111110010101000000101011101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel69[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel69_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel69 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111101010001001010101100011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel69[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel69_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel69 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111101001000011000001010111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel69[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel69_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel69 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111110101011101000100110111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel69[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel69_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel69 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111110110011011110111101000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel69[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel69_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel69 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b10111101001100001101000110111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel69[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel69_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel69 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111110011001111010000100000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel69[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel69_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel69 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111101101010101101001101110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel69[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel69_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel69 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111110001000000101110000101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel69[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel69_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel69 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111110100100110100001100001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel69[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel69_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel69 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111110000111100111011111011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel69[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel69_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel69 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b00111110101011000101010001011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel69[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel69_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel69 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111110101101101011000000111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel69[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel69_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel69 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111110101110101000011010000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel69[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel69_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel69 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111110101010000011100100001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel69[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel69_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel69 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111110011100011001011100011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel69[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel69_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel69 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111110101001110010010011010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel69[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel69_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel69 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b10111101001101011011000010001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel69[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel69_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel69 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111100100110010000110111111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel69[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel69_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel69 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111110010111100100101011110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel69[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel69_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel69 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111110001111000000000111101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel69[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel69_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel69 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111110111101101110101011100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel69[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel69_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel69 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b10111101111000110111111001110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel69[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel69_Valid_Out)
	);
	Adder_64input add_k69(
		.Data1(Data_Out_Kernel69[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel69[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel69[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel69[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel69[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel69[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel69[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel69[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel69[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel69[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel69[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel69[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel69[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel69[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel69[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel69[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel69[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel69[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel69[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel69[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel69[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel69[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel69[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel69[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel69[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel69[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel69[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel69[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel69[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel69[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel69[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel69[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel69[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel69[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel69[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel69[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel69[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel69[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel69[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel69[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel69[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel69[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel69[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel69[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel69[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel69[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel69[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel69[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel69[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel69[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel69[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel69[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel69[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel69[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel69[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel69[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel69[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel69[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel69[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel69[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel69[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel69[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel69[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel69[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel69),
		.Data_Out(add_k69_Data_Out),
		.Valid_Out(add_kernel69_Valid_Out)
	);
	Batch_Norm bn_kernel69(
		.Data_A(32'b00111110011000000011111110100000),
		.Data_B(32'b10111111001101011000000011000101),
		.Data_In(add_k69_Data_Out),
		.Valid_In(add_kernel69_Valid_Out),
		.Data_Out(bn69_Data_Out),
		.Valid_Out(bn69_Valid_Out)
	);
	Relu_Core rl_kernel69(
		.Data_In(bn69_Data_Out),
		.Valid_In(bn69_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*69-1:DATA_WIDHT*68]),
		.Valid_Out(rl69_Valid_Out)
	);
//////////KERNEL70//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel70 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111110111100001101101011100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel70[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel70_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel70 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110011111010011001011001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel70[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel70_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel70 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110100110100101000001011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel70[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel70_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel70 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110100110110111111111011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel70[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel70_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel70 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111101100100011010111010100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel70[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel70_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel70 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110011011010100110010100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel70[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel70_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel70 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111101111010001011000100011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel70[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel70_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel70 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111110001011011101011101000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel70[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel70_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel70 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111101101110111000001101100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel70[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel70_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel70 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111101100111011110100110100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel70[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel70_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel70 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111101100011100111110110010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel70[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel70_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel70 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111110100000101111010101100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel70[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel70_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel70 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111100011000111110100110011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel70[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel70_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel70 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111100000001100001100011100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel70[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel70_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel70 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110101001111100000011101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel70[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel70_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel70 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111101100001111101100110001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel70[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel70_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel70 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111100000000001000110011000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel70[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel70_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel70 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110010010111110111101111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel70[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel70_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel70 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110011011111000011001010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel70[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel70_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel70 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110001101011100001111000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel70[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel70_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel70 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110100111101111110011110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel70[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel70_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel70 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111101101011101101100111011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel70[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel70_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel70 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110111000000110010101110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel70[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel70_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel70 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111101110100100110000100110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel70[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel70_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel70 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111100010101000010101110010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel70[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel70_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel70 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110000110001101101000000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel70[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel70_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel70 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110100100110111111000011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel70[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel70_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel70 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111100111110010111011100011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel70[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel70_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel70 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111110000110100100100111010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel70[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel70_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel70 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111111000000010000100011001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel70[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel70_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel70 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111101011001010101001100100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel70[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel70_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel70 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111101100111101100000100001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel70[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel70_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel70 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b00111101110001001000010101110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel70[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel70_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel70 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b00111110000000010101101011001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel70[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel70_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel70 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111110110011111101000100001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel70[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel70_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel70 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b10111110001101011010110001001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel70[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel70_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel70 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111110000100110000100000101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel70[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel70_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel70 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111101100010110110000000001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel70[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel70_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel70 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b00111101001000111101011000111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel70[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel70_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel70 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b00111100100100010101000011101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel70[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel70_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel70 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111111000110110001101101111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel70[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel70_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel70 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111110010000000110111010011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel70[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel70_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel70 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111101011111000100010110101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel70[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel70_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel70 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111110100100111010111011010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel70[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel70_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel70 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111011111101101100011110001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel70[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel70_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel70 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111110010110001111101000010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel70[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel70_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel70 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111110001011011111101011101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel70[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel70_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel70 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111110100000001100100011111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel70[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel70_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel70 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111101110001001111010011100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel70[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel70_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel70 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111101000110100001001111100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel70[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel70_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel70 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111110100011111101011000100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel70[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel70_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel70 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111100111001100010100100100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel70[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel70_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel70 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111100011100110100001101100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel70[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel70_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel70 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111110010110100001100010001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel70[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel70_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel70 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111110001101011101110101111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel70[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel70_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel70 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b00111001100000111111010011100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel70[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel70_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel70 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111101110110011011110011111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel70[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel70_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel70 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111110000011110010111010001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel70[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel70_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel70 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111101100010101110000100011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel70[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel70_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel70 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111101101111010111111001111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel70[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel70_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel70 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111101101010000111100110001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel70[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel70_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel70 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111101110100010111110110001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel70[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel70_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel70 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111110001010111000010100010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel70[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel70_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel70 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b10111101110110100000100000111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel70[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel70_Valid_Out)
	);
	Adder_64input add_k70(
		.Data1(Data_Out_Kernel70[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel70[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel70[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel70[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel70[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel70[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel70[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel70[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel70[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel70[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel70[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel70[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel70[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel70[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel70[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel70[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel70[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel70[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel70[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel70[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel70[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel70[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel70[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel70[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel70[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel70[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel70[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel70[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel70[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel70[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel70[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel70[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel70[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel70[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel70[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel70[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel70[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel70[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel70[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel70[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel70[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel70[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel70[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel70[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel70[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel70[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel70[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel70[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel70[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel70[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel70[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel70[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel70[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel70[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel70[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel70[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel70[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel70[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel70[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel70[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel70[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel70[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel70[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel70[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel70),
		.Data_Out(add_k70_Data_Out),
		.Valid_Out(add_kernel70_Valid_Out)
	);
	Batch_Norm bn_kernel70(
		.Data_A(32'b00111110100010111011001000001001),
		.Data_B(32'b10111110101001100100001111001100),
		.Data_In(add_k70_Data_Out),
		.Valid_In(add_kernel70_Valid_Out),
		.Data_Out(bn70_Data_Out),
		.Valid_Out(bn70_Valid_Out)
	);
	Relu_Core rl_kernel70(
		.Data_In(bn70_Data_Out),
		.Valid_In(bn70_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*70-1:DATA_WIDHT*69]),
		.Valid_Out(rl70_Valid_Out)
	);
//////////KERNEL71//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel71 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110111010010001110110001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel71[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel71_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel71 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111101101010101001101001001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel71[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel71_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel71 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111001011110111010010101111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel71[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel71_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel71 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111111000011011001110001101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel71[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel71_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel71 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111110010010100111100011100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel71[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel71_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel71 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111101100000010011011000100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel71[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel71_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel71 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111100110101001011111101000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel71[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel71_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel71 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111111000100110101010111001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel71[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel71_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel71 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111111001000001001111000101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel71[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel71_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel71 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111101111100010101000101001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel71[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel71_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel71 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111110100110110010110001111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel71[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel71_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel71 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111110100100101010010101111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel71[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel71_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel71 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110011101110110101000011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel71[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel71_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel71 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111110101010100001110110110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel71[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel71_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel71 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111101100000010011010100010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel71[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel71_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel71 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111110111011111000001111010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel71[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel71_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel71 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111110110011100000110101101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel71[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel71_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel71 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111101001100111111000001111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel71[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel71_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel71 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111001100010100110100011111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel71[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel71_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel71 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111101101011001001111010000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel71[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel71_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel71 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111101111111100011110101110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel71[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel71_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel71 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111110110111001100100011100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel71[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel71_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel71 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111110000000100100101100011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel71[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel71_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel71 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111111010100011011110010111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel71[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel71_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel71 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111110100010001001111011001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel71[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel71_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel71 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111110100101011101101010111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel71[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel71_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel71 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111110010111010000001111100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel71[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel71_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel71 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111111001010110111111011011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel71[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel71_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel71 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111100100011110101001010101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel71[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel71_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel71 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110010101000101010101111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel71[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel71_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel71 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111110010111001011111100011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel71[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel71_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel71 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111110110110001101000011100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel71[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel71_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel71 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111101111110011111011001010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel71[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel71_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel71 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b00111110011011111000100100001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel71[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel71_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel71 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111110110000001100001101100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel71[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel71_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel71 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b10111110011110001001000111010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel71[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel71_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel71 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111101010110001011110010011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel71[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel71_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel71 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111110101011010100101011001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel71[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel71_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel71 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111111010100111001000100100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel71[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel71_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel71 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b00111101111111010010100010101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel71[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel71_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel71 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b10111111011100000111011010010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel71[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel71_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel71 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b10111110111001000100111110100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel71[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel71_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel71 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b00111110101011100010111010101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel71[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel71_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel71 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111110010110100001001100100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel71[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel71_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel71 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b00111110001000001010100000011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel71[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel71_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel71 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b10111110100111111100010111101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel71[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel71_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel71 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111110101001110001011100000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel71[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel71_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel71 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b00111110101010011110010110100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel71[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel71_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel71 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b00111110000000101110101011011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel71[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel71_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel71 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b00111100101010100111011010100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel71[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel71_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel71 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111110011110100110110100101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel71[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel71_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel71 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b10111110101001110110111000100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel71[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel71_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel71 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b00111110000101001001000101111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel71[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel71_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel71 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b00111111000000011100111101100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel71[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel71_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel71 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111110000010011101010001001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel71[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel71_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel71 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b00111110110000000100010010011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel71[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel71_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel71 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b10111110000101010111011011000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel71[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel71_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel71 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b10111110011001000011010111101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel71[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel71_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel71 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b10111110011011110000100111101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel71[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel71_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel71 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b00111110100101001100000111111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel71[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel71_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel71 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111101100001011010001101111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel71[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel71_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel71 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b10111110111011101100101001111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel71[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel71_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel71 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b10111110010111111001100110111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel71[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel71_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel71 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111110010101010001000101100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel71[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel71_Valid_Out)
	);
	Adder_64input add_k71(
		.Data1(Data_Out_Kernel71[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel71[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel71[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel71[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel71[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel71[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel71[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel71[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel71[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel71[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel71[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel71[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel71[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel71[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel71[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel71[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel71[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel71[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel71[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel71[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel71[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel71[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel71[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel71[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel71[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel71[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel71[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel71[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel71[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel71[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel71[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel71[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel71[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel71[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel71[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel71[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel71[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel71[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel71[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel71[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel71[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel71[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel71[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel71[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel71[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel71[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel71[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel71[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel71[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel71[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel71[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel71[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel71[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel71[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel71[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel71[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel71[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel71[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel71[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel71[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel71[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel71[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel71[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel71[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel71),
		.Data_Out(add_k71_Data_Out),
		.Valid_Out(add_kernel71_Valid_Out)
	);
	Batch_Norm bn_kernel71(
		.Data_A(32'b00111110000011101100101101011010),
		.Data_B(32'b00111111011000100000100100111110),
		.Data_In(add_k71_Data_Out),
		.Valid_In(add_kernel71_Valid_Out),
		.Data_Out(bn71_Data_Out),
		.Valid_Out(bn71_Valid_Out)
	);
	Relu_Core rl_kernel71(
		.Data_In(bn71_Data_Out),
		.Valid_In(bn71_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*71-1:DATA_WIDHT*70]),
		.Valid_Out(rl71_Valid_Out)
	);
//////////KERNEL72//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel72 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111101011000000010000101100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel72[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel72_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel72 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111111000100101110100010011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel72[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel72_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel72 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110101101111101001001110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel72[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel72_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel72 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110111111100111110111110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel72[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel72_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel72 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111110000100110011010000110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel72[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel72_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel72 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110000101100000011111001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel72[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel72_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel72 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111110010100100011000100011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel72[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel72_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel72 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111110100101111111010110110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel72[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel72_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel72 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111110100010001101110000011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel72[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel72_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel72 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111101101101000001101000110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel72[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel72_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel72 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111101001101111010111101101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel72[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel72_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel72 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111110011010101110001100111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel72[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel72_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel72 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111101111001010010001110001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel72[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel72_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel72 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111101000010101010001101110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel72[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel72_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel72 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110010001101110000001100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel72[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel72_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel72 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111101110000110110000010011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel72[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel72_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel72 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111110100010101010011111000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel72[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel72_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel72 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111101000111100101101110111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel72[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel72_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel72 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111101111111100101010111011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel72[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel72_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel72 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110001000111000100101010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel72[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel72_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel72 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110001110001110111110111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel72[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel72_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel72 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111101110110011110000101110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel72[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel72_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel72 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111110110100110010110011000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel72[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel72_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel72 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111110111000001010011100111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel72[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel72_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel72 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111010101011001101000101001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel72[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel72_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel72 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111110101000101111101000101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel72[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel72_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel72 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111110111001011001010111010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel72[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel72_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel72 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111110100001111101111110000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel72[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel72_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel72 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111110001000010111101111010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel72[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel72_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel72 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110011101100000010110111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel72[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel72_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel72 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111110101101101111000001101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel72[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel72_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel72 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111110101101100000011010010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel72[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel72_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel72 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111100100001100111001000100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel72[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel72_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel72 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111110010110111111010011010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel72[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel72_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel72 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111110110100100001110011010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel72[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel72_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel72 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111101100100111000001001001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel72[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel72_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel72 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b10111110100001011101001111000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel72[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel72_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel72 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b00111110010001110010010100001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel72[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel72_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel72 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111110111000000111111110101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel72[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel72_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel72 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b00111110010000001100001010111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel72[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel72_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel72 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b10111111010011111010101011100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel72[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel72_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel72 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111110000011101000001111100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel72[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel72_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel72 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b00111101110001101111100111111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel72[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel72_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel72 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b00111100110010110000001100010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel72[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel72_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel72 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b00111110110110100010101011010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel72[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel72_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel72 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b10111110111111101101110011100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel72[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel72_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel72 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b10111101101111000011111011000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel72[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel72_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel72 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b00111110011011001010100011110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel72[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel72_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel72 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111101101000110000011011111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel72[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel72_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel72 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111101010111101100010001001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel72[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel72_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel72 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111101101100100000001101100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel72[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel72_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel72 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b10111110101001010101001010110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel72[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel72_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel72 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111110101111000011111110011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel72[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel72_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel72 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b00111101100001100111110101101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel72[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel72_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel72 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b10111110001010000100110100001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel72[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel72_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel72 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b00111110010000010000101010100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel72[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel72_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel72 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b10111110100011101111011111110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel72[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel72_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel72 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b10111111001000011000011001110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel72[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel72_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel72 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111110100001010101000011000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel72[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel72_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel72 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111110001100101001000001011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel72[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel72_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel72 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b10111101110011111010111011100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel72[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel72_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel72 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111101010111101101111101101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel72[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel72_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel72 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b10111111000000100111010100110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel72[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel72_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel72 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111101000100110010000111000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel72[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel72_Valid_Out)
	);
	Adder_64input add_k72(
		.Data1(Data_Out_Kernel72[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel72[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel72[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel72[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel72[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel72[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel72[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel72[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel72[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel72[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel72[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel72[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel72[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel72[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel72[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel72[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel72[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel72[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel72[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel72[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel72[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel72[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel72[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel72[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel72[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel72[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel72[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel72[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel72[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel72[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel72[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel72[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel72[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel72[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel72[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel72[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel72[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel72[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel72[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel72[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel72[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel72[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel72[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel72[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel72[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel72[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel72[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel72[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel72[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel72[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel72[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel72[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel72[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel72[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel72[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel72[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel72[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel72[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel72[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel72[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel72[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel72[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel72[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel72[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel72),
		.Data_Out(add_k72_Data_Out),
		.Valid_Out(add_kernel72_Valid_Out)
	);
	Batch_Norm bn_kernel72(
		.Data_A(32'b00111110001001101010001011100100),
		.Data_B(32'b00111111001111100110010110000101),
		.Data_In(add_k72_Data_Out),
		.Valid_In(add_kernel72_Valid_Out),
		.Data_Out(bn72_Data_Out),
		.Valid_Out(bn72_Valid_Out)
	);
	Relu_Core rl_kernel72(
		.Data_In(bn72_Data_Out),
		.Valid_In(bn72_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*72-1:DATA_WIDHT*71]),
		.Valid_Out(rl72_Valid_Out)
	);
//////////KERNEL73//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel73 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110010100000000010010011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel73[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel73_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel73 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111101101010100001101101000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel73[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel73_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel73 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111101101001100000101011001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel73[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel73_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel73 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111101100010000010001110110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel73[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel73_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel73 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111110001010010001110001011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel73[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel73_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel73 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110011111001100111110110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel73[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel73_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel73 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111110100111010111101111000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel73[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel73_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel73 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111110100111100011000111100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel73[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel73_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel73 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111101100011100001000011100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel73[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel73_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel73 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110001010110011100110001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel73[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel73_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel73 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111101111110110100111000011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel73[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel73_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel73 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110000000101110101101011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel73[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel73_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel73 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110000111010001111001101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel73[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel73_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel73 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111110101100000111100000110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel73[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel73_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel73 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110110001111100110001010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel73[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel73_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel73 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111111001101100100111001010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel73[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel73_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel73 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111110101100001111010110110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel73[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel73_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel73 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111110100000101111110000100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel73[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel73_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel73 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111101111010011010000100000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel73[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel73_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel73 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110010111111000001001101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel73[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel73_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel73 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110010010010100111100110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel73[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel73_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel73 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111011100010111010001111101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel73[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel73_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel73 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111101011010110001001011111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel73[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel73_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel73 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111111000101011111101100001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel73[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel73_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel73 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111101000110000010110101110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel73[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel73_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel73 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111110100011000110000110010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel73[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel73_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel73 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111111000000101010011110001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel73[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel73_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel73 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111101010110001101101011010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel73[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel73_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel73 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111101100001010111000101000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel73[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel73_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel73 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110100011110100001101100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel73[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel73_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel73 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111110111000100000100000001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel73[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel73_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel73 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111110001011101101101011001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel73[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel73_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel73 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b00111110011000111100001111010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel73[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel73_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel73 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111110110011001101000100010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel73[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel73_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel73 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111111010001111001000100000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel73[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel73_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel73 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111110001011100101111110100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel73[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel73_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel73 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111101100101111111010001000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel73[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel73_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel73 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b00111110100100010011101001100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel73[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel73_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel73 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111110101101000010001101100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel73[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel73_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel73 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b00111110100110111111001111111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel73[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel73_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel73 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b10111110110101011111100001010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel73[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel73_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel73 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111110011001011000101000011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel73[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel73_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel73 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111101011011010010111011100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel73[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel73_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel73 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111110000110110101110011001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel73[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel73_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel73 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b00111111000011100111100101101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel73[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel73_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel73 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b10111110011111010100010011011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel73[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel73_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel73 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b10111110001100011101000000101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel73[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel73_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel73 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b00111110100001111101000010001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel73[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel73_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel73 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111101001000111111111100001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel73[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel73_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel73 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b00111101111100010100101011010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel73[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel73_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel73 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111101110101011000100110011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel73[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel73_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel73 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b10111110101111011111110111110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel73[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel73_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel73 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111110100110001100111010011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel73[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel73_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel73 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b00111110110000010010110010000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel73[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel73_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel73 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b10111101010011111000111000000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel73[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel73_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel73 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b00111110001000101011110011011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel73[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel73_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel73 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b10111111001000001000000110010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel73[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel73_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel73 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b10111110001111101000111000111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel73[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel73_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel73 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111110101110110110010011100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel73[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel73_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel73 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111110000000001010111011111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel73[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel73_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel73 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111110100111011111001100000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel73[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel73_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel73 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111110001100110001011111001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel73[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel73_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel73 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b10111101110100000111111000011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel73[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel73_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel73 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b10111101101101011010101110000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel73[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel73_Valid_Out)
	);
	Adder_64input add_k73(
		.Data1(Data_Out_Kernel73[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel73[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel73[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel73[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel73[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel73[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel73[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel73[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel73[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel73[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel73[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel73[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel73[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel73[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel73[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel73[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel73[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel73[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel73[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel73[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel73[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel73[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel73[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel73[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel73[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel73[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel73[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel73[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel73[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel73[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel73[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel73[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel73[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel73[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel73[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel73[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel73[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel73[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel73[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel73[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel73[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel73[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel73[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel73[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel73[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel73[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel73[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel73[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel73[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel73[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel73[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel73[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel73[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel73[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel73[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel73[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel73[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel73[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel73[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel73[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel73[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel73[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel73[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel73[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel73),
		.Data_Out(add_k73_Data_Out),
		.Valid_Out(add_kernel73_Valid_Out)
	);
	Batch_Norm bn_kernel73(
		.Data_A(32'b00111110001101011001011011010110),
		.Data_B(32'b10111110001001000000111100111011),
		.Data_In(add_k73_Data_Out),
		.Valid_In(add_kernel73_Valid_Out),
		.Data_Out(bn73_Data_Out),
		.Valid_Out(bn73_Valid_Out)
	);
	Relu_Core rl_kernel73(
		.Data_In(bn73_Data_Out),
		.Valid_In(bn73_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*73-1:DATA_WIDHT*72]),
		.Valid_Out(rl73_Valid_Out)
	);
//////////KERNEL74//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel74 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111111001101110001010011011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel74[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel74_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel74 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111110100011010000000111100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel74[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel74_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel74 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110100100100101010000011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel74[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel74_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel74 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111101010011111011011110010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel74[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel74_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel74 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111110000000011001011101110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel74[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel74_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel74 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110100001111100100010100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel74[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel74_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel74 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111110001110011101000111101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel74[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel74_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel74 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111110110100110110001010100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel74[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel74_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel74 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110000111100110011011100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel74[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel74_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel74 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111110001001010110101110001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel74[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel74_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel74 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110100000010000100101001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel74[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel74_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel74 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111101000100000010010011010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel74[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel74_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel74 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111111000000000110111101101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel74[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel74_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel74 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111110011010000010110000111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel74[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel74_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel74 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110100000111011010010000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel74[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel74_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel74 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111110101101011100010011101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel74[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel74_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel74 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110111110011110010000001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel74[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel74_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel74 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110010011100110000000010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel74[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel74_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel74 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111101110111100110101011100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel74[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel74_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel74 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110111001001000001100011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel74[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel74_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel74 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110010111110100000110011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel74[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel74_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel74 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111111001100111100010001010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel74[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel74_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel74 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111011110011001001111001111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel74[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel74_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel74 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111110111000110110110101001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel74[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel74_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel74 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111101111100101101011010000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel74[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel74_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel74 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111110010010101100100010101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel74[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel74_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel74 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111101111101110111100100000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel74[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel74_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel74 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111110001100000101100100100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel74[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel74_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel74 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111101011010001000111101000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel74[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel74_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel74 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111110111101000001110010000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel74[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel74_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel74 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111110010001100101110111000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel74[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel74_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel74 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111101011111000010000111111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel74[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel74_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel74 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b00111110110111110110001111010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel74[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel74_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel74 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111110001001011001010000001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel74[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel74_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel74 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111111001111001100000001100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel74[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel74_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel74 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b10111110110110101000010110110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel74[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel74_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel74 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b10111101111101110100000010101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel74[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel74_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel74 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b00111110110001101001101100111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel74[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel74_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel74 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b00111110010001001011001000001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel74[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel74_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel74 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111110001111010011100010111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel74[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel74_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel74 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111110001011101110101011101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel74[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel74_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel74 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b10111110101111100101100111101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel74[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel74_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel74 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111110001011111111101100011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel74[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel74_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel74 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b00111110000111010110100010111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel74[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel74_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel74 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b00111101101011001100000111110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel74[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel74_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel74 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111111001001111101111010011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel74[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel74_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel74 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111101111001001010111111111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel74[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel74_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel74 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111110100011100101000011001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel74[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel74_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel74 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111110100100101111101101000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel74[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel74_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel74 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111101100100011101110011011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel74[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel74_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel74 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111100100100110000111111101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel74[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel74_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel74 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111110110001011111001100101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel74[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel74_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel74 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b00111110101001010010011110111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel74[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel74_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel74 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b00111110100001100000001000011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel74[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel74_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel74 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111110001111111011010101000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel74[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel74_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel74 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111101100011011110100000101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel74[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel74_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel74 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111111100100000010111010111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel74[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel74_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel74 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111110100110110001100000100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel74[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel74_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel74 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b10111110001111000011111111111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel74[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel74_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel74 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b00111111100000101111000101110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel74[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel74_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel74 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b10111010101110101011000001001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel74[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel74_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel74 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111110001011101001101001001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel74[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel74_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel74 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b10111101101101100110000001100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel74[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel74_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel74 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b10111101010100001100010010100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel74[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel74_Valid_Out)
	);
	Adder_64input add_k74(
		.Data1(Data_Out_Kernel74[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel74[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel74[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel74[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel74[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel74[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel74[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel74[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel74[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel74[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel74[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel74[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel74[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel74[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel74[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel74[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel74[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel74[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel74[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel74[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel74[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel74[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel74[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel74[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel74[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel74[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel74[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel74[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel74[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel74[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel74[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel74[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel74[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel74[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel74[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel74[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel74[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel74[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel74[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel74[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel74[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel74[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel74[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel74[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel74[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel74[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel74[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel74[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel74[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel74[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel74[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel74[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel74[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel74[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel74[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel74[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel74[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel74[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel74[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel74[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel74[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel74[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel74[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel74[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel74),
		.Data_Out(add_k74_Data_Out),
		.Valid_Out(add_kernel74_Valid_Out)
	);
	Batch_Norm bn_kernel74(
		.Data_A(32'b00111110001110010101010101110010),
		.Data_B(32'b10111111101010001010001000011001),
		.Data_In(add_k74_Data_Out),
		.Valid_In(add_kernel74_Valid_Out),
		.Data_Out(bn74_Data_Out),
		.Valid_Out(bn74_Valid_Out)
	);
	Relu_Core rl_kernel74(
		.Data_In(bn74_Data_Out),
		.Valid_In(bn74_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*74-1:DATA_WIDHT*73]),
		.Valid_Out(rl74_Valid_Out)
	);
//////////KERNEL75//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel75 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111111000011001010001010111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel75[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel75_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel75 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110011000101111110101101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel75[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel75_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel75 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110101100011010110111010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel75[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel75_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel75 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111101011001000111100101110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel75[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel75_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel75 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111101001000100001111101001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel75[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel75_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel75 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111100000011001010111110000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel75[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel75_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel75 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111111000100100001100110101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel75[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel75_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel75 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111111001001001100110011111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel75[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel75_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel75 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111110011100000000101011110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel75[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel75_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel75 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110111000110110111100101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel75[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel75_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel75 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110001001110111111011011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel75[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel75_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel75 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110011100011000111010000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel75[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel75_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel75 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111101101011111000000100110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel75[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel75_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel75 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111110110100010100001110000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel75[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel75_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel75 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111101111100010110111000101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel75[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel75_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel75 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111111000000100011111100111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel75[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel75_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel75 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111110101100001101111000100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel75[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel75_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel75 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111011100010100010100111010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel75[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel75_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel75 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111110001111110110101111010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel75[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel75_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel75 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110101101001000100100110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel75[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel75_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel75 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110001100110101100100100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel75[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel75_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel75 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111111000010000001000001010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel75[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel75_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel75 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111110001000011100111111001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel75[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel75_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel75 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111110110110111101101100110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel75[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel75_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel75 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111111100100101010101001001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel75[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel75_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel75 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110101001010010010001000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel75[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel75_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel75 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111110100101011100101101000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel75[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel75_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel75 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111101110101000101110101010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel75[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel75_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel75 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111101101000101101010100001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel75[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel75_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel75 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111111011100000111001010101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel75[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel75_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel75 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111101110011111101010110001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel75[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel75_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel75 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110011100011111111100001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel75[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel75_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel75 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b00111110100001010111000110000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel75[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel75_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel75 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111101101011000001101010011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel75[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel75_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel75 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111110110111111011010011000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel75[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel75_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel75 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b10111101110100101100110110011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel75[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel75_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel75 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b10111110111100010001011011100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel75[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel75_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel75 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111111000010011011011001011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel75[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel75_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel75 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111110111100010001101001111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel75[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel75_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel75 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b00111101110110100100010101101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel75[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel75_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel75 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b10111110100000111110010001000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel75[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel75_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel75 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b10111101111000000011010110110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel75[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel75_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel75 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111011110111111101100010110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel75[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel75_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel75 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111110110001001011010101100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel75[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel75_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel75 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b00111101101100111110011001110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel75[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel75_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel75 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b10111110101111000000100000100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel75[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel75_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel75 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b10111101011000110100111101010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel75[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel75_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel75 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b00111110011111100110110010010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel75[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel75_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel75 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b00111110101010011000010010011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel75[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel75_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel75 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b00111110101000010001001000111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel75[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel75_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel75 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b10111110000110110111110001100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel75[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel75_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel75 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b10111110101000101100110101000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel75[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel75_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel75 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111110010011000000010111110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel75[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel75_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel75 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b00111110010110100011010101000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel75[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel75_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel75 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111011110010001110111100111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel75[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel75_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel75 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b00111110011001100011101100010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel75[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel75_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel75 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b10111111001100011111001010100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel75[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel75_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel75 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b10111110101110000111010111111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel75[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel75_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel75 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111011010101011010000111110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel75[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel75_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel75 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111101110010010111100000011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel75[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel75_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel75 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b10111101001110111101101110101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel75[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel75_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel75 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111110001100100111101011001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel75[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel75_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel75 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111110001110000010110110001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel75[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel75_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel75 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b10111110010100111011010001100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel75[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel75_Valid_Out)
	);
	Adder_64input add_k75(
		.Data1(Data_Out_Kernel75[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel75[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel75[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel75[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel75[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel75[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel75[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel75[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel75[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel75[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel75[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel75[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel75[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel75[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel75[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel75[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel75[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel75[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel75[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel75[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel75[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel75[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel75[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel75[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel75[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel75[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel75[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel75[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel75[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel75[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel75[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel75[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel75[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel75[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel75[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel75[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel75[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel75[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel75[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel75[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel75[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel75[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel75[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel75[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel75[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel75[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel75[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel75[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel75[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel75[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel75[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel75[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel75[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel75[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel75[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel75[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel75[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel75[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel75[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel75[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel75[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel75[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel75[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel75[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel75),
		.Data_Out(add_k75_Data_Out),
		.Valid_Out(add_kernel75_Valid_Out)
	);
	Batch_Norm bn_kernel75(
		.Data_A(32'b00111110000010010001011100101010),
		.Data_B(32'b00111110101011010000001110001111),
		.Data_In(add_k75_Data_Out),
		.Valid_In(add_kernel75_Valid_Out),
		.Data_Out(bn75_Data_Out),
		.Valid_Out(bn75_Valid_Out)
	);
	Relu_Core rl_kernel75(
		.Data_In(bn75_Data_Out),
		.Valid_In(bn75_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*75-1:DATA_WIDHT*74]),
		.Valid_Out(rl75_Valid_Out)
	);
//////////KERNEL76//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel76 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111110101110111110111001010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel76[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel76_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel76 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110000100111100001111111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel76[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel76_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel76 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111101110011110010110011001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel76[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel76_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel76 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110001000011110000001100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel76[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel76_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel76 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111101111010110111001011010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel76[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel76_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel76 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111100110100010100000011111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel76[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel76_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel76 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111110001011001001110000000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel76[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel76_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel76 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111110010010001001111010110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel76[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel76_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel76 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111101110010111111100100010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel76[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel76_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel76 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111110010010000111101100001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel76[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel76_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel76 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111101100110000011010011010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel76[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel76_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel76 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111100100001110110111011000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel76[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel76_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel76 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111100111110010001001011110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel76[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel76_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel76 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111110001100110111101111010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel76[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel76_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel76 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111010101100010010101100111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel76[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel76_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel76 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111110100011110100010010101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel76[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel76_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel76 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110000111100011110001100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel76[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel76_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel76 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111101101110101010000111001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel76[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel76_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel76 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111101001010110000100100111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel76[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel76_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel76 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111101100101110010011011011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel76[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel76_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel76 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110101010011101111011001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel76[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel76_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel76 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111101100111011001001011011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel76[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel76_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel76 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110100011110010011011100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel76[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel76_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel76 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111101110010011110001110010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel76[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel76_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel76 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111100110011111110001111100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel76[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel76_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel76 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110101100001010000010111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel76[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel76_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel76 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111111000100001011010100110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel76[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel76_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel76 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111101110000001111100010001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel76[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel76_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel76 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111110001000010011110000110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel76[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel76_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel76 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111101010011001010111001001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel76[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel76_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel76 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111111000000111010010101100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel76[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel76_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel76 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110101010010111001110010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel76[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel76_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel76 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111110000101101110001011000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel76[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel76_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel76 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b00111110101001100011011011000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel76[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel76_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel76 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111110111101101111011000111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel76[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel76_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel76 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b10111101111110001110010100001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel76[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel76_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel76 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111110100011101000000010111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel76[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel76_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel76 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111110001111110101100010111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel76[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel76_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel76 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b00111110000111101111001011110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel76[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel76_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel76 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111110000010110100101000010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel76[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel76_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel76 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111111000111110100101000111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel76[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel76_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel76 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111101101001011111001110101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel76[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel76_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel76 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111101010010001011010100100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel76[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel76_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel76 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111100110010010001000010110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel76[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel76_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel76 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111110010100010110111010111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel76[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel76_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel76 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111110101010010000110111111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel76[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel76_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel76 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111110001101111011000000011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel76[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel76_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel76 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111110001101110000111001000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel76[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel76_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel76 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b00111101011000001100010110100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel76[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel76_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel76 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b00111101000110011100001100000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel76[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel76_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel76 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111101111011011010001101101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel76[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel76_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel76 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111110010101111110010011010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel76[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel76_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel76 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b00111110100011000001010101011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel76[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel76_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel76 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111110111110111001000000110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel76[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel76_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel76 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111110010000111100000001111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel76[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel76_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel76 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111110001001111001110010010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel76[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel76_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel76 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111110110010001000000000111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel76[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel76_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel76 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111110010101000011110010101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel76[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel76_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel76 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b10111110011001000111010011000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel76[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel76_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel76 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b00111110001110100111101000101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel76[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel76_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel76 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111110001010011110100000010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel76[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel76_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel76 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111110000100000001000001100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel76[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel76_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel76 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111110101111111000001000000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel76[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel76_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel76 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111101011110110100101101010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel76[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel76_Valid_Out)
	);
	Adder_64input add_k76(
		.Data1(Data_Out_Kernel76[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel76[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel76[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel76[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel76[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel76[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel76[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel76[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel76[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel76[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel76[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel76[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel76[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel76[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel76[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel76[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel76[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel76[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel76[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel76[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel76[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel76[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel76[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel76[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel76[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel76[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel76[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel76[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel76[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel76[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel76[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel76[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel76[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel76[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel76[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel76[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel76[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel76[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel76[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel76[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel76[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel76[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel76[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel76[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel76[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel76[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel76[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel76[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel76[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel76[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel76[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel76[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel76[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel76[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel76[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel76[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel76[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel76[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel76[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel76[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel76[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel76[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel76[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel76[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel76),
		.Data_Out(add_k76_Data_Out),
		.Valid_Out(add_kernel76_Valid_Out)
	);
	Batch_Norm bn_kernel76(
		.Data_A(32'b00111110010101000000100101101100),
		.Data_B(32'b10111111001111000110000110010010),
		.Data_In(add_k76_Data_Out),
		.Valid_In(add_kernel76_Valid_Out),
		.Data_Out(bn76_Data_Out),
		.Valid_Out(bn76_Valid_Out)
	);
	Relu_Core rl_kernel76(
		.Data_In(bn76_Data_Out),
		.Valid_In(bn76_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*76-1:DATA_WIDHT*75]),
		.Valid_Out(rl76_Valid_Out)
	);
//////////KERNEL77//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel77 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111110100110110101001001110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel77[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel77_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel77 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110100011111110011001001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel77[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel77_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel77 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110110011011101101010001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel77[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel77_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel77 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110110101101001110111000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel77[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel77_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel77 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111101100110100001010100110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel77[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel77_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel77 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111101111010011110011000110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel77[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel77_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel77 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111101100000000111100110111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel77[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel77_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel77 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111100001001011101101111101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel77[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel77_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel77 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111101110001111101101111000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel77[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel77_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel77 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111101110101011100111100010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel77[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel77_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel77 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111101000101010011010110001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel77[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel77_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel77 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111101100111100110010000111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel77[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel77_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel77 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111100101001010000101000001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel77[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel77_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel77 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111101001001101111101010100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel77[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel77_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel77 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110100000001000101111100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel77[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel77_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel77 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111101000110001101111000011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel77[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel77_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel77 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110000010110010010111100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel77[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel77_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel77 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110001000011000100000111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel77[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel77_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel77 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111101011111101110010111000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel77[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel77_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel77 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110001101000101001100001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel77[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel77_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel77 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110111000000101110101000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel77[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel77_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel77 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111101100010111110010010001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel77[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel77_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel77 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110101111000001111100100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel77[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel77_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel77 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111110010100111111010011010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel77[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel77_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel77 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111100110001110011001111111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel77[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel77_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel77 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110100111010000001101000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel77[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel77_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel77 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110111001011111111100010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel77[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel77_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel77 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110100000111010101001001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel77[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel77_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel77 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111110001111010010111111010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel77[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel77_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel77 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111110100010011010101010100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel77[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel77_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel77 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111110010001101100111011111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel77[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel77_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel77 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110110000011010100011001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel77[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel77_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel77 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111110101100001101101000110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel77[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel77_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel77 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b00111110010011011001000111000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel77[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel77_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel77 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111111000011100100001010001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel77[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel77_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel77 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b10111110100110101110000111101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel77[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel77_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel77 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111110001101011100110111101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel77[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel77_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel77 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111101110101010101111001000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel77[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel77_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel77 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b00111110001111001000010001000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel77[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel77_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel77 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111101100110100000111011010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel77[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel77_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel77 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111111001001111111111010111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel77[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel77_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel77 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111110100101000110000001000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel77[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel77_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel77 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b00111101000010111101001111011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel77[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel77_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel77 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111101110000100110011001110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel77[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel77_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel77 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111110111001000100011110101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel77[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel77_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel77 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111110101000000101001100010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel77[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel77_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel77 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b10111101111111110111101110111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel77[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel77_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel77 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111110101011110110100100101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel77[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel77_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel77 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111110001000000110110110101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel77[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel77_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel77 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b00111101010000100100010110100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel77[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel77_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel77 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111110101100111001000110110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel77[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel77_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel77 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111110001011111001011110101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel77[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel77_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel77 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b00111110100011010100010100100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel77[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel77_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel77 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111111000000010110110110100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel77[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel77_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel77 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111110000111010011111000101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel77[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel77_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel77 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111110101000110000010111101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel77[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel77_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel77 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111110100010011001001000010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel77[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel77_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel77 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111110000110010111110111111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel77[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel77_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel77 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111110000100110011000100100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel77[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel77_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel77 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b00111101001010000101011100010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel77[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel77_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel77 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111110100011011110101101101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel77[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel77_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel77 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b10111101100010010111000111011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel77[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel77_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel77 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111101110000011100001000011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel77[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel77_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel77 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b10111101111110101111001001000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel77[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel77_Valid_Out)
	);
	Adder_64input add_k77(
		.Data1(Data_Out_Kernel77[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel77[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel77[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel77[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel77[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel77[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel77[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel77[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel77[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel77[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel77[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel77[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel77[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel77[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel77[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel77[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel77[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel77[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel77[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel77[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel77[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel77[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel77[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel77[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel77[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel77[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel77[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel77[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel77[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel77[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel77[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel77[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel77[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel77[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel77[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel77[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel77[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel77[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel77[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel77[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel77[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel77[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel77[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel77[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel77[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel77[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel77[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel77[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel77[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel77[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel77[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel77[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel77[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel77[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel77[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel77[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel77[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel77[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel77[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel77[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel77[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel77[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel77[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel77[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel77),
		.Data_Out(add_k77_Data_Out),
		.Valid_Out(add_kernel77_Valid_Out)
	);
	Batch_Norm bn_kernel77(
		.Data_A(32'b00111110010000110001010100001110),
		.Data_B(32'b10111111000010101001010011100111),
		.Data_In(add_k77_Data_Out),
		.Valid_In(add_kernel77_Valid_Out),
		.Data_Out(bn77_Data_Out),
		.Valid_Out(bn77_Valid_Out)
	);
	Relu_Core rl_kernel77(
		.Data_In(bn77_Data_Out),
		.Valid_In(bn77_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*77-1:DATA_WIDHT*76]),
		.Valid_Out(rl77_Valid_Out)
	);
//////////KERNEL78//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel78 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110011010100001110110001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel78[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel78_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel78 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111101110101011100110111111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel78[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel78_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel78 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110010111010110111011001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel78[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel78_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel78 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111100100010101101010001110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel78[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel78_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel78 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111101001110010100011011011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel78[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel78_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel78 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111100000111000100101111010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel78[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel78_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel78 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111111001000010111010011101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel78[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel78_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel78 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111101100101100101110000000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel78[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel78_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel78 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111110111100010111101000011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel78[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel78_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel78 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110110000101110010110111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel78[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel78_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel78 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111111100110100110011001011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel78[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel78_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel78 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111110110101011111000011100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel78[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel78_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel78 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111101101010100001010001011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel78[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel78_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel78 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111111001011110010111010111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel78[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel78_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel78 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110100010010001101011001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel78[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel78_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel78 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111101100000101010000010101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel78[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel78_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel78 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111111000010110010100011110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel78[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel78_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel78 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111110110000100111001100110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel78[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel78_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel78 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110110100000100010000111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel78[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel78_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel78 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111110010011001011010110010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel78[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel78_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel78 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110110001001111011110100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel78[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel78_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel78 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111110101011111010000101110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel78[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel78_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel78 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111101100100010111111000010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel78[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel78_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel78 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111111001101000000110100001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel78[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel78_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel78 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111101001001110111111010011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel78[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel78_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel78 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111110100100010010110000001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel78[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel78_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel78 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111111000110100001101010010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel78[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel78_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel78 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111101011100111000000010011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel78[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel78_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel78 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111110000001011110101100101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel78[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel78_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel78 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111101100010000110110111110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel78[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel78_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel78 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111101101101101110000011111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel78[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel78_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel78 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111110100001101011100011111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel78[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel78_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel78 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b00111101000011011100101001101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel78[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel78_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel78 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111110001101011011011111101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel78[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel78_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel78 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111101010011111001111100000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel78[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel78_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel78 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111101000101101101001001011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel78[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel78_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel78 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111101001111011100100011111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel78[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel78_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel78 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111101111010011100101000010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel78[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel78_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel78 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111110110101101000001011101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel78[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel78_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel78 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b00111110110010100010001111011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel78[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel78_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel78 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b10111111100001100101110011100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel78[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel78_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel78 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b10111110111100111000000000000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel78[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel78_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel78 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b00111110000011010011110110011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel78[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel78_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel78 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111110001110110101101000100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel78[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel78_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel78 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b00111101000011010000111001100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel78[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel78_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel78 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b10111110001101000100000111001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel78[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel78_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel78 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111110001110110000100100101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel78[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel78_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel78 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b00111111000111000011011101011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel78[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel78_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel78 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111110000111001100100101101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel78[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel78_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel78 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b00111110011011111010111010001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel78[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel78_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel78 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b10111101111110011000011101011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel78[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel78_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel78 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111101110010000001111100110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel78[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel78_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel78 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b00111110001100101001011010101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel78[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel78_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel78 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b00111110101110101000010111100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel78[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel78_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel78 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b10111111000011000000101110111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel78[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel78_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel78 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111110011000010010101100011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel78[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel78_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel78 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111101101000011110011000101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel78[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel78_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel78 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b10111110011001001100001110100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel78[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel78_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel78 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111101111000000011100000100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel78[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel78_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel78 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111110100000110101111100111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel78[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel78_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel78 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b10111110000001010101111111010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel78[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel78_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel78 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b10111110100000010010101111110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel78[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel78_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel78 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b10111110101100000100110101011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel78[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel78_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel78 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111110110101001011111111101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel78[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel78_Valid_Out)
	);
	Adder_64input add_k78(
		.Data1(Data_Out_Kernel78[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel78[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel78[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel78[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel78[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel78[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel78[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel78[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel78[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel78[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel78[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel78[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel78[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel78[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel78[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel78[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel78[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel78[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel78[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel78[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel78[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel78[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel78[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel78[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel78[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel78[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel78[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel78[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel78[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel78[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel78[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel78[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel78[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel78[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel78[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel78[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel78[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel78[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel78[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel78[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel78[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel78[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel78[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel78[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel78[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel78[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel78[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel78[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel78[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel78[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel78[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel78[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel78[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel78[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel78[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel78[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel78[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel78[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel78[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel78[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel78[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel78[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel78[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel78[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel78),
		.Data_Out(add_k78_Data_Out),
		.Valid_Out(add_kernel78_Valid_Out)
	);
	Batch_Norm bn_kernel78(
		.Data_A(32'b00111110000111111101110101000111),
		.Data_B(32'b00111111100010101010010101000100),
		.Data_In(add_k78_Data_Out),
		.Valid_In(add_kernel78_Valid_Out),
		.Data_Out(bn78_Data_Out),
		.Valid_Out(bn78_Valid_Out)
	);
	Relu_Core rl_kernel78(
		.Data_In(bn78_Data_Out),
		.Valid_In(bn78_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*78-1:DATA_WIDHT*77]),
		.Valid_Out(rl78_Valid_Out)
	);
//////////KERNEL79//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel79 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111101010110001011111101110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel79[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel79_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel79 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110100000101111111101011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel79[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel79_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel79 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110110001111100101101101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel79[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel79_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel79 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110101100000101111110010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel79[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel79_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel79 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111110011101001110101010001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel79[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel79_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel79 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110001101100001111010111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel79[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel79_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel79 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111111000100111001000111100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel79[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel79_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel79 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111101011111010011010000100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel79[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel79_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel79 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111111010110110101001001101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel79[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel79_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel79 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110001110100101010001001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel79[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel79_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel79 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110101000110010001000001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel79[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel79_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel79 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111110100111011101000000101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel79[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel79_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel79 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110000010010100011010001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel79[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel79_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel79 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111100101011001101010101101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel79[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel79_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel79 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111101001101100110100100100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel79[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel79_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel79 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111110011011101101101000010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel79[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel79_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel79 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111111000111101110011010100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel79[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel79_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel79 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111110000100000001011101111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel79[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel79_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel79 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111101100101110110111001110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel79[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel79_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel79 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111100111000010111101100000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel79[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel79_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel79 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111111001000100100011011000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel79[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel79_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel79 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111110000111101101111011001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel79[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel79_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel79 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111111000010011000100000010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel79[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel79_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel79 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111111100111101010011101001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel79[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel79_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel79 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111101101111010011001001111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel79[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel79_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel79 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111101111000011101101010100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel79[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel79_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel79 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110101011101101111100010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel79[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel79_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel79 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110001001011110001111010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel79[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel79_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel79 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111110010111100110001011000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel79[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel79_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel79 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110011001110110011111000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel79[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel79_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel79 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111110100101001101001011101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel79[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel79_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel79 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111101110011111111000000001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel79[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel79_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel79 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111110101101110110001010110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel79[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel79_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel79 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b00111110110110101000010101100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel79[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel79_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel79 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111110000001100001000111111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel79[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel79_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel79 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111100011111000101011011101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel79[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel79_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel79 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111111000111000110001011000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel79[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel79_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel79 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111110011011001001010110001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel79[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel79_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel79 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b00111110000100000011101001110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel79[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel79_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel79 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b00111101100001111011100110001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel79[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel79_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel79 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111111001111010011100011001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel79[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel79_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel79 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b10111110000111101110000010000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel79[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel79_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel79 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111110001100111110000100111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel79[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel79_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel79 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111101010011011110001010111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel79[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel79_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel79 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111110111100101010111110000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel79[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel79_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel79 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111110110100011110110010000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel79[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel79_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel79 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111101010001110000001101101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel79[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel79_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel79 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111110100111101010011101100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel79[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel79_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel79 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111110101010111000010110111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel79[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel79_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel79 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111110001010010100000010000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel79[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel79_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel79 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111101011101011101010111001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel79[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel79_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel79 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111110100000001001011010100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel79[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel79_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel79 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111101100110100011100101010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel79[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel79_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel79 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111111001001111000101011001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel79[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel79_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel79 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111100010101001011010111100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel79[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel79_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel79 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111110111101011001100100001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel79[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel79_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel79 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111110011111000101111011101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel79[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel79_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel79 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111110010010010010101111010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel79[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel79_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel79 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b10111100100110001100011110010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel79[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel79_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel79 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b00111110101000100000001000110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel79[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel79_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel79 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b10111110000101010110111011011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel79[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel79_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel79 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111100111100110100001100110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel79[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel79_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel79 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111101101001101100001011101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel79[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel79_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel79 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111110000010100111000101101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel79[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel79_Valid_Out)
	);
	Adder_64input add_k79(
		.Data1(Data_Out_Kernel79[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel79[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel79[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel79[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel79[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel79[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel79[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel79[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel79[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel79[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel79[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel79[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel79[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel79[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel79[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel79[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel79[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel79[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel79[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel79[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel79[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel79[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel79[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel79[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel79[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel79[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel79[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel79[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel79[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel79[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel79[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel79[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel79[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel79[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel79[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel79[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel79[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel79[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel79[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel79[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel79[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel79[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel79[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel79[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel79[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel79[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel79[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel79[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel79[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel79[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel79[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel79[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel79[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel79[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel79[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel79[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel79[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel79[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel79[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel79[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel79[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel79[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel79[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel79[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel79),
		.Data_Out(add_k79_Data_Out),
		.Valid_Out(add_kernel79_Valid_Out)
	);
	Batch_Norm bn_kernel79(
		.Data_A(32'b00111101111001100001000100011010),
		.Data_B(32'b00111100110101010100001010011000),
		.Data_In(add_k79_Data_Out),
		.Valid_In(add_kernel79_Valid_Out),
		.Data_Out(bn79_Data_Out),
		.Valid_Out(bn79_Valid_Out)
	);
	Relu_Core rl_kernel79(
		.Data_In(bn79_Data_Out),
		.Valid_In(bn79_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*79-1:DATA_WIDHT*78]),
		.Valid_Out(rl79_Valid_Out)
	);
//////////KERNEL80//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel80 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110101111000101001111000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel80[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel80_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel80 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111101111010111111001100100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel80[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel80_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel80 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111100101011110000010111001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel80[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel80_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel80 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110101000110111001011111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel80[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel80_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel80 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111011110000011100000111110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel80[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel80_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel80 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111101101100111000000000110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel80[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel80_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel80 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111110001011001101101100011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel80[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel80_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel80 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111101010100110100000010000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel80[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel80_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel80 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111111000101101000100000010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel80[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel80_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel80 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111101000101001101011101101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel80[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel80_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel80 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110001011010111101001011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel80[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel80_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel80 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110000101110110100000000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel80[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel80_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel80 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111101010111000111101011110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel80[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel80_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel80 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111110100100101000110101010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel80[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel80_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel80 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110010100001011101011001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel80[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel80_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel80 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111110000000001011111101010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel80[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel80_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel80 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111111000110100000000100111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel80[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel80_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel80 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111100101100010011011100100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel80[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel80_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel80 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111110100001001010100011010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel80[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel80_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel80 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111101100100000011011101011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel80[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel80_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel80 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110100110000110110110000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel80[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel80_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel80 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111101100111100110100110110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel80[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel80_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel80 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111110010100111011000101010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel80[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel80_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel80 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111110100001101100000010101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel80[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel80_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel80 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111110100011100100010000110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel80[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel80_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel80 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111110011101101010101001101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel80[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel80_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel80 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111110100000000011010101011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel80[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel80_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel80 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111110100101011011001111111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel80[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel80_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel80 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111100011111011011100110101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel80[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel80_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel80 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110100001101011111001010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel80[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel80_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel80 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111110000111010111100001010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel80[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel80_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel80 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111001110011100011000001111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel80[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel80_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel80 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b00111110110011001001101010001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel80[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel80_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel80 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111110100000000011110100111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel80[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel80_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel80 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111111000110100011010100011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel80[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel80_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel80 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111110000010000001100010001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel80[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel80_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel80 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b10111110100101101011001100000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel80[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel80_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel80 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b00111100010010110100100011001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel80[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel80_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel80 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111111000001011000010100010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel80[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel80_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel80 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b00111101011111100100000110111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel80[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel80_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel80 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b10111110100001000111100111110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel80[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel80_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel80 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111101110010111101110111110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel80[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel80_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel80 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b00111110010100111100000001101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel80[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel80_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel80 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111101110111111110111000001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel80[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel80_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel80 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b00111110101111011010000110111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel80[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel80_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel80 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b10111101111011100110110110100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel80[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel80_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel80 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b10111110100000101110100110001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel80[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel80_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel80 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b00111110111011011001110010001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel80[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel80_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel80 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111011100000101101110000101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel80[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel80_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel80 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b00111110001001100000010101010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel80[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel80_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel80 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111110001010010100101100011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel80[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel80_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel80 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b10111110101001101000010111111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel80[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel80_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel80 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111101101000111000011010111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel80[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel80_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel80 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b00111110100001110000100101111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel80[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel80_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel80 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111100111001110100100101100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel80[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel80_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel80 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b00111101111000111111110101110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel80[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel80_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel80 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b10111110111100001110111100000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel80[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel80_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel80 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b10111110110010010000011011101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel80[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel80_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel80 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111110111011011001110000001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel80[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel80_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel80 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111101011010110011011101001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel80[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel80_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel80 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b10111011100110000110101010000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel80[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel80_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel80 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111110010011000110000000001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel80[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel80_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel80 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111101011101101101010001101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel80[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel80_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel80 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111100000100010100001101111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel80[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel80_Valid_Out)
	);
	Adder_64input add_k80(
		.Data1(Data_Out_Kernel80[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel80[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel80[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel80[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel80[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel80[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel80[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel80[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel80[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel80[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel80[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel80[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel80[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel80[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel80[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel80[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel80[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel80[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel80[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel80[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel80[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel80[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel80[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel80[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel80[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel80[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel80[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel80[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel80[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel80[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel80[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel80[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel80[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel80[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel80[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel80[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel80[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel80[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel80[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel80[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel80[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel80[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel80[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel80[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel80[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel80[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel80[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel80[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel80[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel80[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel80[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel80[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel80[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel80[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel80[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel80[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel80[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel80[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel80[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel80[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel80[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel80[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel80[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel80[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel80),
		.Data_Out(add_k80_Data_Out),
		.Valid_Out(add_kernel80_Valid_Out)
	);
	Batch_Norm bn_kernel80(
		.Data_A(32'b00111110001111100101011101100110),
		.Data_B(32'b10111110001100000001100101000110),
		.Data_In(add_k80_Data_Out),
		.Valid_In(add_kernel80_Valid_Out),
		.Data_Out(bn80_Data_Out),
		.Valid_Out(bn80_Valid_Out)
	);
	Relu_Core rl_kernel80(
		.Data_In(bn80_Data_Out),
		.Valid_In(bn80_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*80-1:DATA_WIDHT*79]),
		.Valid_Out(rl80_Valid_Out)
	);
//////////KERNEL81//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel81 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110101000000110101100100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel81[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel81_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel81 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111110001001101110101110101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel81[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel81_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel81 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110101001011100001010110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel81[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel81_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel81 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110010001010001110010100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel81[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel81_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel81 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111101010000110100110000000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel81[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel81_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel81 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111101110011011001100100101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel81[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel81_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel81 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111110010101000110101111100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel81[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel81_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel81 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111101101100100110001011110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel81[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel81_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel81 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111110000110100110101000011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel81[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel81_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel81 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110100110101011111000100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel81[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel81_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel81 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110001011010010010010101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel81[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel81_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel81 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111101101111011110001101101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel81[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel81_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel81 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111101111100001111111111001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel81[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel81_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel81 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111110011011111001000110001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel81[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel81_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel81 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110010010011001010100111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel81[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel81_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel81 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111110110000101110100100001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel81[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel81_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel81 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111110110001010000111100110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel81[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel81_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel81 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111101100110011101011001111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel81[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel81_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel81 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111010010010001011101011001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel81[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel81_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel81 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111101100000101001101111111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel81[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel81_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel81 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110111011101011010000000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel81[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel81_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel81 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111110010101001110000010110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel81[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel81_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel81 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111110011101111110101001010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel81[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel81_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel81 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111110111000010110111001001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel81[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel81_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel81 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111110100001001111100110000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel81[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel81_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel81 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111110010010000101100001101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel81[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel81_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel81 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111110111001010011001100001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel81[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel81_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel81 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111110110101010010110000100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel81[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel81_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel81 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111110001011010011111101100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel81[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel81_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel81 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110101000011001100110001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel81[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel81_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel81 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111101101101011110011001011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel81[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel81_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel81 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111110000111110010100111000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel81[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel81_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel81 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b00111110100000010000010011111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel81[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel81_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel81 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111110101110101011000111011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel81[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel81_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel81 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111111010100011110100001001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel81[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel81_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel81 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111110001110000000010101110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel81[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel81_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel81 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b10111110001001010101101011011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel81[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel81_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel81 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111110000001011111011111001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel81[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel81_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel81 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111110110001101101001010011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel81[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel81_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel81 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b00111110011100010000011111100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel81[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel81_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel81 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b10111110110000010111000100100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel81[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel81_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel81 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111110010010110010001100011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel81[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel81_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel81 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111100111001110100001001110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel81[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel81_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel81 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111110001000111011001001000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel81[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel81_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel81 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b00111110100110111111110101100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel81[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel81_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel81 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b10111110100111100010011101110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel81[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel81_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel81 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b10111101111100011000111010000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel81[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel81_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel81 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b00111110101011100101101100100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel81[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel81_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel81 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b00111101110011110000011101000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel81[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel81_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel81 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b00111110011010011010010001110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel81[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel81_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel81 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111101110110101000001110001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel81[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel81_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel81 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b10111110110101001000010010101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel81[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel81_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel81 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111110100010010001101011100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel81[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel81_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel81 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b00111110100111011101110111000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel81[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel81_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel81 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111011101101000101101111011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel81[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel81_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel81 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b00111101111111010111100011111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel81[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel81_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel81 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b10111111000011110110011010000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel81[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel81_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel81 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b10111110100001000101111101000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel81[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel81_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel81 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111110101011011111010011110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel81[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel81_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel81 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111011111100110111110000110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel81[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel81_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel81 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111101111111011111011100011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel81[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel81_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel81 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111101110101010001010101111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel81[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel81_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel81 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111101011111100000110001001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel81[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel81_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel81 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111110000001001111011111010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel81[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel81_Valid_Out)
	);
	Adder_64input add_k81(
		.Data1(Data_Out_Kernel81[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel81[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel81[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel81[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel81[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel81[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel81[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel81[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel81[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel81[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel81[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel81[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel81[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel81[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel81[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel81[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel81[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel81[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel81[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel81[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel81[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel81[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel81[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel81[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel81[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel81[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel81[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel81[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel81[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel81[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel81[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel81[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel81[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel81[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel81[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel81[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel81[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel81[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel81[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel81[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel81[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel81[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel81[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel81[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel81[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel81[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel81[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel81[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel81[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel81[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel81[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel81[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel81[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel81[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel81[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel81[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel81[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel81[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel81[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel81[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel81[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel81[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel81[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel81[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel81),
		.Data_Out(add_k81_Data_Out),
		.Valid_Out(add_kernel81_Valid_Out)
	);
	Batch_Norm bn_kernel81(
		.Data_A(32'b00111110001001110110000011000000),
		.Data_B(32'b00111110100111110001111100001010),
		.Data_In(add_k81_Data_Out),
		.Valid_In(add_kernel81_Valid_Out),
		.Data_Out(bn81_Data_Out),
		.Valid_Out(bn81_Valid_Out)
	);
	Relu_Core rl_kernel81(
		.Data_In(bn81_Data_Out),
		.Valid_In(bn81_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*81-1:DATA_WIDHT*80]),
		.Valid_Out(rl81_Valid_Out)
	);
//////////KERNEL82//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel82 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111110100111101010001000010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel82[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel82_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel82 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110101110011100100101111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel82[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel82_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel82 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110001100001110011010101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel82[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel82_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel82 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110011011001111011101111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel82[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel82_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel82 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111101010101010110100001000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel82[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel82_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel82 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111101010110000110001001000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel82[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel82_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel82 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111110010000111000001001100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel82[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel82_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel82 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111101000011100110101101110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel82[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel82_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel82 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110111010111101001000110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel82[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel82_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel82 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111100100010110110011100110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel82[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel82_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel82 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110011101011010110100000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel82[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel82_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel82 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111100100011110100001110000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel82[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel82_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel82 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110000011000001101011010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel82[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel82_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel82 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111101011000011100111010001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel82[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel82_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel82 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111101111101111100101000001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel82[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel82_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel82 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111101111110100101111000101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel82[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel82_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel82 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110100011001111110000100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel82[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel82_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel82 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111110011011010011110110101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel82[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel82_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel82 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111110010010101101010000010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel82[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel82_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel82 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110111010110001111000100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel82[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel82_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel82 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110110101111000001111100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel82[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel82_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel82 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111110100010010011000011011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel82[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel82_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel82 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111101111010010000011110101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel82[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel82_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel82 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111110111010011001011110000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel82[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel82_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel82 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111110011111111010000000111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel82[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel82_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel82 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110011111100111010101001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel82[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel82_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel82 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111111000000000010011001110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel82[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel82_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel82 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110110001111100000101101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel82[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel82_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel82 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111100011011111011100100010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel82[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel82_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel82 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111101001100011010111000011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel82[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel82_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel82 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111110010000011010000010110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel82[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel82_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel82 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110000111000111110100011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel82[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel82_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel82 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111111000111111010001011000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel82[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel82_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel82 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b00111111000110110100110000000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel82[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel82_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel82 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111111001010010011100010110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel82[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel82_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel82 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111101111111010101110101011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel82[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel82_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel82 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111110100110100011100011111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel82[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel82_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel82 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111101111101111100100100110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel82[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel82_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel82 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b00111101100000011111000011110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel82[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel82_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel82 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b00111110000000101111010110111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel82[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel82_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel82 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111110111100001001110011111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel82[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel82_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel82 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111101111011100111010111011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel82[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel82_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel82 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b00111101001001101100000001100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel82[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel82_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel82 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b00111101010011001111011000011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel82[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel82_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel82 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111111000110110011010100000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel82[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel82_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel82 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111110111110011101011110101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel82[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel82_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel82 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111110100001100000001101010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel82[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel82_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel82 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111111001001101001100011100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel82[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel82_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel82 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111110000001110101101011010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel82[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel82_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel82 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111011111101111000111101000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel82[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel82_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel82 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b10111101001000111010100001101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel82[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel82_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel82 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111111000101001011010010001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel82[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel82_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel82 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b00111110001111111010101110000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel82[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel82_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel82 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111110111101100101001000101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel82[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel82_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel82 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b10111110000101111100011010000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel82[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel82_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel82 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111110101110101010100100101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel82[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel82_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel82 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111110100000010011010101111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel82[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel82_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel82 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b10111100110000001110110010000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel82[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel82_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel82 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b10111110010000011111100001001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel82[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel82_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel82 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b00111110000111010011000011111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel82[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel82_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel82 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b10111100011011111111100011000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel82[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel82_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel82 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111101010010100111001111100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel82[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel82_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel82 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b10111100011001100101000010111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel82[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel82_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel82 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111100011010101011011011110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel82[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel82_Valid_Out)
	);
	Adder_64input add_k82(
		.Data1(Data_Out_Kernel82[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel82[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel82[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel82[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel82[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel82[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel82[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel82[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel82[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel82[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel82[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel82[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel82[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel82[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel82[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel82[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel82[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel82[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel82[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel82[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel82[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel82[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel82[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel82[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel82[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel82[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel82[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel82[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel82[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel82[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel82[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel82[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel82[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel82[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel82[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel82[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel82[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel82[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel82[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel82[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel82[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel82[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel82[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel82[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel82[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel82[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel82[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel82[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel82[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel82[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel82[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel82[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel82[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel82[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel82[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel82[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel82[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel82[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel82[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel82[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel82[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel82[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel82[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel82[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel82),
		.Data_Out(add_k82_Data_Out),
		.Valid_Out(add_kernel82_Valid_Out)
	);
	Batch_Norm bn_kernel82(
		.Data_A(32'b00111110001010010111111001101111),
		.Data_B(32'b10111110101100110111010111110010),
		.Data_In(add_k82_Data_Out),
		.Valid_In(add_kernel82_Valid_Out),
		.Data_Out(bn82_Data_Out),
		.Valid_Out(bn82_Valid_Out)
	);
	Relu_Core rl_kernel82(
		.Data_In(bn82_Data_Out),
		.Valid_In(bn82_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*82-1:DATA_WIDHT*81]),
		.Valid_Out(rl82_Valid_Out)
	);
//////////KERNEL83//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel83 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111111000011011011111001110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel83[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel83_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel83 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110001011011111100101000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel83[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel83_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel83 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110000100111011011101101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel83[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel83_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel83 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110101110101001010011010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel83[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel83_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel83 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111110000101111111101001010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel83[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel83_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel83 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110000111110111010011001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel83[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel83_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel83 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111101100100000001100110110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel83[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel83_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel83 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111101011011010010101011001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel83[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel83_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel83 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110011010101011000011011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel83[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel83_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel83 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110010110101110111011000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel83[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel83_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel83 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111101011001011001010000111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel83[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel83_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel83 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111110010100011110111110011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel83[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel83_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel83 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110011110111111111001110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel83[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel83_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel83 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111101001110111100111011011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel83[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel83_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel83 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110100011010111100100101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel83[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel83_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel83 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111100010000011001110110000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel83[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel83_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel83 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110111110011010101010001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel83[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel83_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel83 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110000100011101011100100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel83[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel83_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel83 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110001100100100011101110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel83[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel83_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel83 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110010100110110101000001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel83[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel83_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel83 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110000111110001111011110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel83[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel83_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel83 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111101110111010000111101001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel83[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel83_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel83 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110111101110111111101111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel83[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel83_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel83 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111101111001111110100101111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel83[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel83_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel83 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111110100101111110001101101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel83[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel83_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel83 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110010001010110000111110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel83[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel83_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel83 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110001110100111011110000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel83[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel83_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel83 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111101110010100001101110010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel83[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel83_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel83 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111110011011011111001110011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel83[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel83_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel83 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111110011010111010101011000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel83[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel83_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel83 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111101110111101110001111110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel83[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel83_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel83 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111101011001101011110100110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel83[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel83_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel83 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b00111011111110110001101001100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel83[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel83_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel83 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b00111101000000111001011011100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel83[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel83_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel83 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111110110010100001111111000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel83[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel83_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel83 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b10111101100011101000100111111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel83[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel83_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel83 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111110110100110011010100001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel83[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel83_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel83 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111100000111010111101111011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel83[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel83_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel83 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b00111101111101001001110110100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel83[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel83_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel83 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111110000010011000111100101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel83[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel83_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel83 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111111000111110011010010110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel83[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel83_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel83 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111110011100111101001000111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel83[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel83_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel83 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111110001001101101010011010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel83[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel83_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel83 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111110001010110100011101101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel83[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel83_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel83 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111101100001011101000111110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel83[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel83_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel83 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111101011110010110010110001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel83[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel83_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel83 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111110110100111001010001010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel83[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel83_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel83 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111110000001000110101011001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel83[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel83_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel83 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111110000110011010110110111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel83[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel83_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel83 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111101100110111011011100110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel83[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel83_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel83 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111110010011000001100010010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel83[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel83_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel83 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b10111101000100011000010101100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel83[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel83_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel83 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111101111100111001101110010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel83[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel83_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel83 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111110011010111000010010001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel83[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel83_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel83 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111110000100100111001100100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel83[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel83_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel83 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b00111110001110011010000011101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel83[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel83_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel83 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111110100010101011001011001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel83[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel83_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel83 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111110001101101100111110000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel83[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel83_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel83 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111100101011011000011100011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel83[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel83_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel83 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b00111101011011001000100111111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel83[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel83_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel83 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111110010111101000101110001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel83[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel83_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel83 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111101100111010111011110001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel83[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel83_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel83 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111110001001101011101001111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel83[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel83_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel83 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b10111101011100100011100111010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel83[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel83_Valid_Out)
	);
	Adder_64input add_k83(
		.Data1(Data_Out_Kernel83[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel83[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel83[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel83[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel83[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel83[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel83[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel83[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel83[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel83[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel83[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel83[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel83[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel83[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel83[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel83[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel83[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel83[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel83[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel83[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel83[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel83[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel83[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel83[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel83[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel83[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel83[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel83[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel83[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel83[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel83[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel83[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel83[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel83[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel83[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel83[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel83[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel83[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel83[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel83[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel83[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel83[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel83[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel83[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel83[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel83[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel83[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel83[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel83[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel83[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel83[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel83[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel83[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel83[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel83[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel83[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel83[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel83[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel83[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel83[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel83[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel83[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel83[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel83[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel83),
		.Data_Out(add_k83_Data_Out),
		.Valid_Out(add_kernel83_Valid_Out)
	);
	Batch_Norm bn_kernel83(
		.Data_A(32'b00111110011000110100001101100011),
		.Data_B(32'b10111111001101100111011011111011),
		.Data_In(add_k83_Data_Out),
		.Valid_In(add_kernel83_Valid_Out),
		.Data_Out(bn83_Data_Out),
		.Valid_Out(bn83_Valid_Out)
	);
	Relu_Core rl_kernel83(
		.Data_In(bn83_Data_Out),
		.Valid_In(bn83_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*83-1:DATA_WIDHT*82]),
		.Valid_Out(rl83_Valid_Out)
	);
//////////KERNEL84//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel84 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111110100010110110111010111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel84[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel84_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel84 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110010111000001000110011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel84[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel84_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel84 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111101111001010110100000110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel84[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel84_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel84 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111101111110100011011010111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel84[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel84_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel84 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111110001011101001111111011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel84[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel84_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel84 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111100000011010010101011010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel84[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel84_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel84 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111110000111011011001101111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel84[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel84_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel84 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111011101000001110011101001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel84[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel84_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel84 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111101100010000100111110011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel84[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel84_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel84 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111110101001101010111100111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel84[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel84_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel84 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111101000010010001101101001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel84[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel84_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel84 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111100111010010011101000011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel84[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel84_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel84 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111101100111100110110010001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel84[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel84_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel84 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111101011001110101000100000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel84[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel84_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel84 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110100110001111011011011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel84[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel84_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel84 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111110001001110001101000100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel84[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel84_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel84 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111101101100001001011011001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel84[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel84_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel84 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111101111010011011000101011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel84[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel84_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel84 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110011011000011100010010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel84[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel84_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel84 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111101101110000111010100111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel84[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel84_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel84 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110100101010010001000101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel84[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel84_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel84 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111101101001011000111001111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel84[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel84_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel84 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110011001010111000101111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel84[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel84_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel84 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111110011110110111010001110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel84[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel84_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel84 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111101010101111010101100111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel84[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel84_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel84 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110100111100100010111111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel84[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel84_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel84 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110111000001110011110100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel84[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel84_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel84 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111101101110101000111111111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel84[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel84_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel84 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111101011100010111111010111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel84[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel84_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel84 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111110101110011001100111000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel84[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel84_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel84 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111110100100110100011110010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel84[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel84_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel84 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110100111101110010100010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel84[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel84_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel84 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111101001001011100010000101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel84[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel84_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel84 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b00111110010010110111111000101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel84[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel84_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel84 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111110101001011111001001001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel84[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel84_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel84 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b10111101111101100111011111000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel84[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel84_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel84 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111101100100101001011100111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel84[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel84_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel84 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111101001011001110100011011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel84[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel84_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel84 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b00111101101100100111010111110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel84[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel84_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel84 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b00111101101001100101001110000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel84[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel84_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel84 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111111001100010101010011000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel84[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel84_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel84 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111101100111101101111010011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel84[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel84_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel84 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b00111010101110110010111010010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel84[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel84_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel84 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111101101110101010110001001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel84[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel84_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel84 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111110100001001010101111000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel84[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel84_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel84 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111110111011001110010100111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel84[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel84_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel84 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111110001011010111011011101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel84[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel84_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel84 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111110011000101010111111001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel84[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel84_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel84 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b00111101101100001100111101100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel84[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel84_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel84 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111101011010000111101000000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel84[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel84_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel84 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111110001001101001111000011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel84[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel84_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel84 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111110011101110101001100010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel84[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel84_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel84 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b00111110010100011101101011001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel84[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel84_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel84 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111110111111001100101110111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel84[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel84_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel84 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111101101000110101111101011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel84[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel84_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel84 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111110010100010101001001010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel84[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel84_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel84 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111110101000000110100001011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel84[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel84_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel84 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111101111010100011101100100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel84[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel84_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel84 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b10111110010110000001100101111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel84[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel84_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel84 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111101000010100101101001111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel84[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel84_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel84 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111110000100110010011010010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel84[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel84_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel84 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111100101000110111110101111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel84[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel84_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel84 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111110110111010110001011011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel84[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel84_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel84 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b10111101100110011000111111101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel84[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel84_Valid_Out)
	);
	Adder_64input add_k84(
		.Data1(Data_Out_Kernel84[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel84[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel84[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel84[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel84[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel84[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel84[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel84[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel84[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel84[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel84[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel84[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel84[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel84[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel84[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel84[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel84[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel84[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel84[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel84[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel84[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel84[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel84[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel84[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel84[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel84[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel84[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel84[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel84[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel84[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel84[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel84[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel84[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel84[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel84[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel84[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel84[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel84[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel84[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel84[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel84[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel84[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel84[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel84[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel84[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel84[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel84[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel84[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel84[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel84[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel84[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel84[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel84[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel84[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel84[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel84[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel84[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel84[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel84[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel84[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel84[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel84[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel84[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel84[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel84),
		.Data_Out(add_k84_Data_Out),
		.Valid_Out(add_kernel84_Valid_Out)
	);
	Batch_Norm bn_kernel84(
		.Data_A(32'b00111110010111110010000001101011),
		.Data_B(32'b10111110110011011100000100011011),
		.Data_In(add_k84_Data_Out),
		.Valid_In(add_kernel84_Valid_Out),
		.Data_Out(bn84_Data_Out),
		.Valid_Out(bn84_Valid_Out)
	);
	Relu_Core rl_kernel84(
		.Data_In(bn84_Data_Out),
		.Valid_In(bn84_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*84-1:DATA_WIDHT*83]),
		.Valid_Out(rl84_Valid_Out)
	);
//////////KERNEL85//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel85 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111110101011110001010100011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel85[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel85_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel85 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110100101010010000100011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel85[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel85_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel85 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111101011100111110001100100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel85[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel85_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel85 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111111000011001110011101110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel85[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel85_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel85 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111110000100101001101111100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel85[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel85_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel85 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111101111110011011001011100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel85[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel85_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel85 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111101011011010110101100110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel85[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel85_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel85 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111110000000100001100001000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel85[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel85_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel85 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111101110110101111110101111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel85[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel85_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel85 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111101100110110100110000001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel85[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel85_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel85 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110011010000110101110001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel85[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel85_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel85 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110101100100110011011110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel85[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel85_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel85 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111101000101000001110011100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel85[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel85_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel85 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111110101001011000101000010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel85[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel85_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel85 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110001000110101110001011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel85[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel85_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel85 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111101111110001101000111011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel85[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel85_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel85 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111111000110011100000110110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel85[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel85_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel85 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111110000001111100101101101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel85[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel85_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel85 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111101011001110010000000010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel85[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel85_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel85 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110011111111100101100110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel85[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel85_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel85 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110110011100101001110001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel85[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel85_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel85 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111110000011001111011011001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel85[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel85_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel85 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110001000100111011100001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel85[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel85_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel85 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111110011000011110100010111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel85[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel85_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel85 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111110010110100001100001010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel85[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel85_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel85 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110101010101001000111100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel85[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel85_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel85 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111101100111010010100010011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel85[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel85_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel85 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111110001111100010010110011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel85[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel85_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel85 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111110011010010001101001100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel85[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel85_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel85 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111101111110111010011001000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel85[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel85_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel85 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111101110110011010000101000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel85[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel85_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel85 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111111000110110100011000101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel85[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel85_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel85 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111110110100011111010001000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel85[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel85_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel85 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b00111101101011010011111010111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel85[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel85_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel85 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111110100111000101000010000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel85[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel85_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel85 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111110000011011010001010011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel85[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel85_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel85 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111110001100011111110011111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel85[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel85_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel85 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111101010010100000110100111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel85[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel85_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel85 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b00111110110011101111000100010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel85[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel85_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel85 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b00111011111111101011111001110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel85[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel85_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel85 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111111001001000101111011101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel85[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel85_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel85 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111111000111110111000111010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel85[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel85_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel85 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111101000000100000111010111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel85[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel85_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel85 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b00111110000011111001101010110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel85[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel85_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel85 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111111000101111011000110000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel85[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel85_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel85 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111110100101111001111100011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel85[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel85_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel85 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111110000110100101001101111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel85[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel85_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel85 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111110110011011011001100000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel85[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel85_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel85 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111101011011101101100100000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel85[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel85_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel85 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b00111100000001011010000011111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel85[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel85_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel85 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111110010011011100111000011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel85[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel85_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel85 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111110101011011001111010001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel85[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel85_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel85 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111101000101000010110100110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel85[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel85_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel85 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111110111110011111111100111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel85[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel85_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel85 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b10111101000001010001101000111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel85[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel85_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel85 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111110001010011101100001010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel85[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel85_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel85 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111110011010101111101010110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel85[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel85_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel85 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111101100101110111000001101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel85[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel85_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel85 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111101110110111000001101000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel85[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel85_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel85 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111110001111011001011001010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel85[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel85_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel85 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111110001001001100110110101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel85[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel85_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel85 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b10111100010011101110110100110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel85[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel85_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel85 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111110100010001000001110101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel85[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel85_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel85 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b10111110011000001010111110101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel85[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel85_Valid_Out)
	);
	Adder_64input add_k85(
		.Data1(Data_Out_Kernel85[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel85[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel85[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel85[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel85[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel85[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel85[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel85[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel85[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel85[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel85[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel85[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel85[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel85[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel85[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel85[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel85[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel85[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel85[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel85[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel85[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel85[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel85[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel85[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel85[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel85[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel85[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel85[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel85[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel85[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel85[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel85[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel85[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel85[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel85[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel85[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel85[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel85[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel85[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel85[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel85[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel85[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel85[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel85[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel85[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel85[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel85[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel85[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel85[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel85[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel85[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel85[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel85[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel85[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel85[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel85[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel85[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel85[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel85[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel85[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel85[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel85[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel85[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel85[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel85),
		.Data_Out(add_k85_Data_Out),
		.Valid_Out(add_kernel85_Valid_Out)
	);
	Batch_Norm bn_kernel85(
		.Data_A(32'b00111110001100111000000001110010),
		.Data_B(32'b10111111010101111100110100110110),
		.Data_In(add_k85_Data_Out),
		.Valid_In(add_kernel85_Valid_Out),
		.Data_Out(bn85_Data_Out),
		.Valid_Out(bn85_Valid_Out)
	);
	Relu_Core rl_kernel85(
		.Data_In(bn85_Data_Out),
		.Valid_In(bn85_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*85-1:DATA_WIDHT*84]),
		.Valid_Out(rl85_Valid_Out)
	);
//////////KERNEL86//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel86 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110110111011010111000110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel86[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel86_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel86 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111110110111100101000010010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel86[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel86_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel86 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110100111011010001011001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel86[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel86_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel86 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110110111100101010111000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel86[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel86_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel86 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111110000110001101000100011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel86[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel86_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel86 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111101101100010001010101100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel86[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel86_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel86 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111110001010001010011110001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel86[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel86_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel86 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111101010000101010010000001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel86[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel86_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel86 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111110101001000110000010010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel86[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel86_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel86 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110010101010100010100110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel86[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel86_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel86 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111100011100111010101010111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel86[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel86_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel86 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110001110011110010010101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel86[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel86_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel86 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111101100100101000101100111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel86[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel86_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel86 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111100110111000000011110001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel86[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel86_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel86 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111111000000001010001101110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel86[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel86_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel86 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111101001010101111011010101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel86[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel86_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel86 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111110110100010000010100100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel86[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel86_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel86 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111101100000000100011100010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel86[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel86_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel86 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111100010101100001000100010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel86[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel86_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel86 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111101010101100010111110101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel86[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel86_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel86 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110101010101010011001111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel86[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel86_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel86 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111100110110010011001111010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel86[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel86_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel86 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111110101011100000101101011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel86[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel86_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel86 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111101101010100001111100100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel86[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel86_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel86 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111110010100010001011101000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel86[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel86_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel86 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111110010000110100101111011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel86[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel86_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel86 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111110101011111010100111101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel86[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel86_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel86 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111110101011011011000001010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel86[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel86_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel86 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111110000111010100100101101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel86[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel86_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel86 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110000101000001001011011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel86[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel86_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel86 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111101000011111111000000111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel86[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel86_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel86 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111110100111001001000111110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel86[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel86_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel86 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b00111110011111111000010000010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel86[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel86_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel86 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111110011110100101100001111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel86[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel86_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel86 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111110101100111111111001000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel86[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel86_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel86 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111101110100010111100010011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel86[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel86_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel86 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b10111110100110101011101010000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel86[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel86_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel86 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111110000001011011010101111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel86[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel86_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel86 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111110010011001011100010011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel86[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel86_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel86 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111011101011110010111001110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel86[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel86_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel86 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b10111110111111101011010110100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel86[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel86_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel86 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b10111110010110101001111101110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel86[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel86_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel86 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b00111101011011010111101100001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel86[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel86_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel86 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111100110011011111011011000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel86[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel86_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel86 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b00111110011001001100011010011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel86[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel86_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel86 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b10111110010001000111011001111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel86[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel86_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel86 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b10111110011000010111010001100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel86[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel86_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel86 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b00111110100000110001111100010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel86[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel86_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel86 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111100001010011010001111011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel86[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel86_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel86 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111101100011101011100001010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel86[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel86_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel86 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111101000110011011111101101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel86[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel86_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel86 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b10111110011010100100100000000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel86[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel86_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel86 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111110010101111010001010111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel86[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel86_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel86 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b00111101110011000101000000011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel86[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel86_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel86 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b10111101000010001010001001010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel86[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel86_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel86 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111101100100101011001111011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel86[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel86_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel86 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b10111110100101100001001011100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel86[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel86_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel86 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b10111110110101110001001101100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel86[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel86_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel86 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111101111111001110111111001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel86[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel86_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel86 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111101011111101011110011110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel86[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel86_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel86 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b10111101111011110100001110011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel86[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel86_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel86 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111101000110010011111001111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel86[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel86_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel86 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111101101111100100000110010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel86[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel86_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel86 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111110100001101011101011101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel86[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel86_Valid_Out)
	);
	Adder_64input add_k86(
		.Data1(Data_Out_Kernel86[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel86[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel86[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel86[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel86[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel86[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel86[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel86[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel86[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel86[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel86[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel86[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel86[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel86[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel86[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel86[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel86[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel86[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel86[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel86[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel86[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel86[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel86[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel86[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel86[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel86[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel86[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel86[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel86[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel86[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel86[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel86[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel86[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel86[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel86[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel86[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel86[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel86[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel86[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel86[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel86[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel86[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel86[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel86[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel86[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel86[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel86[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel86[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel86[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel86[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel86[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel86[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel86[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel86[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel86[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel86[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel86[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel86[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel86[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel86[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel86[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel86[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel86[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel86[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel86),
		.Data_Out(add_k86_Data_Out),
		.Valid_Out(add_kernel86_Valid_Out)
	);
	Batch_Norm bn_kernel86(
		.Data_A(32'b00111110010100001111001100001010),
		.Data_B(32'b00111111000100000010101010111110),
		.Data_In(add_k86_Data_Out),
		.Valid_In(add_kernel86_Valid_Out),
		.Data_Out(bn86_Data_Out),
		.Valid_Out(bn86_Valid_Out)
	);
	Relu_Core rl_kernel86(
		.Data_In(bn86_Data_Out),
		.Valid_In(bn86_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*86-1:DATA_WIDHT*85]),
		.Valid_Out(rl86_Valid_Out)
	);
//////////KERNEL87//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel87 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111110101110111010111010011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel87[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel87_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel87 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110011001000101111101111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel87[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel87_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel87 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110010101001010110010110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel87[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel87_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel87 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110111010111010110100110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel87[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel87_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel87 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111101111010010100011111111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel87[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel87_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel87 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110100101110101010001011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel87[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel87_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel87 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111101100101001101100100111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel87[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel87_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel87 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111110000111001001010011101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel87[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel87_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel87 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111101100011010011010110000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel87[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel87_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel87 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111101100011110010000111101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel87[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel87_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel87 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110011000101000100000001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel87[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel87_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel87 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111100001100111011111100100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel87[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel87_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel87 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111100001000100011100000000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel87[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel87_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel87 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111100110011001000000111000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel87[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel87_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel87 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110100110111110111100010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel87[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel87_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel87 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111101110110010100010001010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel87[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel87_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel87 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110100110100111001010110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel87[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel87_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel87 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110001001101011111100011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel87[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel87_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel87 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110000010010011010111011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel87[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel87_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel87 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110100000111101011000100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel87[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel87_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel87 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110100000001000101010101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel87[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel87_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel87 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111101111111101001111010000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel87[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel87_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel87 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110110101000111101000110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel87[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel87_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel87 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111101110110101010100010011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel87[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel87_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel87 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111101011010101100011010001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel87[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel87_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel87 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110000101010000001111100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel87[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel87_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel87 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110010001101000111010110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel87[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel87_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel87 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111101001111100101110010100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel87[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel87_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel87 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111101101111110010101001110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel87[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel87_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel87 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111111000000100100001010101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel87[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel87_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel87 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111110010011101110100100011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel87[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel87_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel87 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110010011110100110111010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel87[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel87_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel87 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111101100100000000010011011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel87[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel87_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel87 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b00111100100101011001010111111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel87[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel87_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel87 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111110110010111011110111110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel87[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel87_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel87 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b10111110001011101000001000011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel87[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel87_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel87 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111101111110001101001011101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel87[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel87_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel87 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b00111101101101010100000101100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel87[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel87_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel87 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b00111110100111110011111101011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel87[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel87_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel87 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b00111010101011001101110000011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel87[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel87_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel87 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111111001000110110110010110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel87[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel87_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel87 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111110100001011010011000011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel87[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel87_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel87 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111101110000011100011011010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel87[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel87_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel87 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111101110011000010110001000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel87[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel87_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel87 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111110010110100100100100000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel87[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel87_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel87 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111110000111010110110001101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel87[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel87_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel87 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111101110001010001000100100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel87[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel87_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel87 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111110100100111000100000100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel87[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel87_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel87 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111110010111111111111010110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel87[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel87_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel87 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111101100000010001010100011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel87[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel87_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel87 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111110100101110110101100101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel87[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel87_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel87 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111101101011001001010000100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel87[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel87_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel87 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b00111101001001111111011000000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel87[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel87_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel87 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111110100110111001100100000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel87[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel87_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel87 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111110100101001011110001001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel87[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel87_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel87 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111101010001000000000000101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel87[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel87_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel87 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111101110001110000110000011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel87[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel87_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel87 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111110000000101100101101100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel87[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel87_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel87 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111110100101100000110011110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel87[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel87_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel87 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111101101110011010010000001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel87[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel87_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel87 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111110010101101000011111111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel87[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel87_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel87 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111110001110110001001010010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel87[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel87_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel87 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111110101010011101011110000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel87[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel87_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel87 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b10111110000011001000001000101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel87[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel87_Valid_Out)
	);
	Adder_64input add_k87(
		.Data1(Data_Out_Kernel87[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel87[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel87[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel87[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel87[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel87[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel87[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel87[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel87[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel87[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel87[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel87[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel87[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel87[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel87[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel87[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel87[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel87[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel87[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel87[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel87[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel87[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel87[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel87[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel87[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel87[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel87[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel87[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel87[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel87[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel87[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel87[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel87[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel87[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel87[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel87[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel87[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel87[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel87[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel87[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel87[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel87[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel87[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel87[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel87[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel87[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel87[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel87[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel87[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel87[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel87[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel87[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel87[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel87[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel87[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel87[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel87[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel87[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel87[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel87[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel87[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel87[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel87[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel87[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel87),
		.Data_Out(add_k87_Data_Out),
		.Valid_Out(add_kernel87_Valid_Out)
	);
	Batch_Norm bn_kernel87(
		.Data_A(32'b00111110011000111110111100100000),
		.Data_B(32'b10111111010000111001010101010100),
		.Data_In(add_k87_Data_Out),
		.Valid_In(add_kernel87_Valid_Out),
		.Data_Out(bn87_Data_Out),
		.Valid_Out(bn87_Valid_Out)
	);
	Relu_Core rl_kernel87(
		.Data_In(bn87_Data_Out),
		.Valid_In(bn87_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*87-1:DATA_WIDHT*86]),
		.Valid_Out(rl87_Valid_Out)
	);
//////////KERNEL88//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel88 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111101000011000101001011111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel88[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel88_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel88 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111110001111010111111111111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel88[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel88_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel88 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111101101110000100000110001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel88[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel88_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel88 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110100101100110111001000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel88[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel88_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel88 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111110100110101011011111101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel88[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel88_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel88 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111101011000001010011110001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel88[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel88_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel88 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111110101101101111000010010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel88[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel88_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel88 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111101101100111001110111111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel88[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel88_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel88 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110101010101000101011101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel88[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel88_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel88 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111111001100001010101110001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel88[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel88_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel88 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111111011110101110001000111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel88[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel88_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel88 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110101111101100001010111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel88[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel88_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel88 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110010011110110011101011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel88[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel88_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel88 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111110001100001001010011110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel88[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel88_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel88 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111101100111111010101001000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel88[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel88_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel88 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111100110100111111000010001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel88[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel88_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel88 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111110100000100111011000101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel88[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel88_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel88 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111101001101111001001110110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel88[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel88_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel88 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111111010101000101010110000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel88[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel88_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel88 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111101111111110110110110111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel88[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel88_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel88 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110000010101000000001011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel88[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel88_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel88 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111110001111011101110000110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel88[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel88_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel88 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111101111000100001100101100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel88[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel88_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel88 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111101000101101000100101011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel88[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel88_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel88 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111110101010000111101001100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel88[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel88_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel88 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111011111111011010111000011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel88[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel88_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel88 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111110110100100110100001100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel88[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel88_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel88 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111100111000111100000111001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel88[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel88_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel88 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111111001000000111000001010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel88[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel88_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel88 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110111101000010111100001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel88[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel88_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel88 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111110110101011011111011001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel88[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel88_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel88 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111111010010001000101101110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel88[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel88_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel88 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111101111100110001011100000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel88[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel88_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel88 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111111001011010010100000111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel88[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel88_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel88 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111110101011011111001101000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel88[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel88_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel88 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111110100111001010101110100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel88[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel88_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel88 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b10111110111111101000001100000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel88[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel88_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel88 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111110010000000011110010001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel88[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel88_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel88 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111110101000010100100010101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel88[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel88_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel88 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b00111110101010001010010110100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel88[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel88_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel88 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b10111101110011011011000110111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel88[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel88_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel88 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b10111110001011100100100001001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel88[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel88_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel88 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111110000010110000001110000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel88[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel88_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel88 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111101110011111111110001000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel88[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel88_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel88 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b00111110101000011000011100101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel88[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel88_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel88 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b10111110001111011111000001100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel88[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel88_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel88 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b10111110010000101011001001110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel88[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel88_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel88 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b00111110110001110011010101110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel88[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel88_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel88 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b00111110001001010011110101100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel88[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel88_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel88 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111110111110101110100110111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel88[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel88_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel88 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b10111110110000011010011000110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel88[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel88_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel88 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b10111110001011100011110001101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel88[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel88_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel88 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111111010001001111110011001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel88[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel88_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel88 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111110101011010101000010111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel88[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel88_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel88 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111101111011101011100100011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel88[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel88_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel88 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b00111101111000110001010110111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel88[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel88_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel88 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111100101000100011101010101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel88[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel88_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel88 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111110110011110111110111101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel88[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel88_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel88 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b10111101110100101101011100000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel88[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel88_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel88 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b00111110101100100111111000011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel88[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel88_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel88 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111110001110001010100010110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel88[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel88_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel88 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b10111110010100010110100011100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel88[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel88_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel88 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b10111110101010101110110100101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel88[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel88_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel88 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b10111110111110000101100010110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel88[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel88_Valid_Out)
	);
	Adder_64input add_k88(
		.Data1(Data_Out_Kernel88[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel88[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel88[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel88[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel88[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel88[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel88[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel88[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel88[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel88[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel88[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel88[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel88[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel88[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel88[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel88[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel88[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel88[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel88[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel88[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel88[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel88[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel88[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel88[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel88[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel88[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel88[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel88[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel88[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel88[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel88[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel88[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel88[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel88[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel88[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel88[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel88[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel88[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel88[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel88[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel88[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel88[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel88[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel88[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel88[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel88[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel88[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel88[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel88[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel88[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel88[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel88[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel88[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel88[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel88[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel88[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel88[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel88[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel88[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel88[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel88[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel88[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel88[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel88[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel88),
		.Data_Out(add_k88_Data_Out),
		.Valid_Out(add_kernel88_Valid_Out)
	);
	Batch_Norm bn_kernel88(
		.Data_A(32'b00111110010010110100101011100011),
		.Data_B(32'b00111111100001101000110000110101),
		.Data_In(add_k88_Data_Out),
		.Valid_In(add_kernel88_Valid_Out),
		.Data_Out(bn88_Data_Out),
		.Valid_Out(bn88_Valid_Out)
	);
	Relu_Core rl_kernel88(
		.Data_In(bn88_Data_Out),
		.Valid_In(bn88_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*88-1:DATA_WIDHT*87]),
		.Valid_Out(rl88_Valid_Out)
	);
//////////KERNEL89//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel89 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110010001001000010100000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel89[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel89_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel89 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111101101101100010000011100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel89[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel89_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel89 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110100001110011111101101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel89[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel89_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel89 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110000101001011001100101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel89[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel89_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel89 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111100111011001110111111100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel89[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel89_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel89 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111100001010110001000101101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel89[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel89_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel89 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111101001101101001011110000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel89[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel89_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel89 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111110010101111000001111101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel89[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel89_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel89 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111110011101001101110111111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel89[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel89_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel89 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110101110110011011000111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel89[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel89_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel89 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111111010000111100100110110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel89[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel89_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel89 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111110011101100000100011001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel89[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel89_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel89 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111101110101001101000010100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel89[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel89_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel89 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111101001001000011111111001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel89[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel89_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel89 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110000100101110011101010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel89[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel89_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel89 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111110100000100010110000001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel89[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel89_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel89 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111111000101010111110100111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel89[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel89_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel89 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111110001011010010101000010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel89[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel89_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel89 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111111000111001000000001000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel89[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel89_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel89 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111110000101110001101001000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel89[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel89_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel89 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110011000100101000101100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel89[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel89_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel89 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111110100111011011011101111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel89[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel89_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel89 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111101011011011111000011101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel89[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel89_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel89 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111110111110010001100111111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel89[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel89_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel89 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111001111110000000011010010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel89[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel89_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel89 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111110101000100001111010111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel89[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel89_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel89 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111111010000001111001100010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel89[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel89_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel89 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110101110001011011110101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel89[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel89_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel89 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111110101011010010001001010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel89[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel89_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel89 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110111000001110110000110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel89[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel89_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel89 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111101000101111001011110101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel89[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel89_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel89 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111111010011010001000100110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel89[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel89_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel89 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111101001111110000000010010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel89[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel89_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel89 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111101010011011001010100001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel89[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel89_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel89 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111111000101011101010010100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel89[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel89_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel89 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111100100111100101100001010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel89[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel89_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel89 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b10111110000010000011011001100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel89[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel89_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel89 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111110110110100011110010011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel89[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel89_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel89 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111111010100100111110011010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel89[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel89_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel89 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b00111110110001101010100010011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel89[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel89_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel89 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b10111111011010001100110010011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel89[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel89_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel89 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b10111111010001010010000101111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel89[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel89_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel89 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b00111110001001000110000111011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel89[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel89_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel89 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111101101011010100100010100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel89[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel89_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel89 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b00111110101000100101110100100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel89[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel89_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel89 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b10111110001001111111101011111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel89[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel89_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel89 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111110010011011110001111011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel89[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel89_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel89 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b00111111000110100110101101000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel89[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel89_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel89 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b00111110010000110100100010011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel89[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel89_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel89 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111110100100101111101001100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel89[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel89_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel89 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111100101111101011101010111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel89[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel89_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel89 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b10111101110000101111010100110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel89[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel89_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel89 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111100100000001001110100101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel89[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel89_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel89 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b00111110010100100110101010101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel89[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel89_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel89 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111101110111110110010011010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel89[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel89_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel89 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b00111101111110100110100001000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel89[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel89_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel89 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b10111100101010010000101011001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel89[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel89_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel89 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111011110001111000001110001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel89[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel89_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel89 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b10111110011000111011111010001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel89[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel89_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel89 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b00111110101000110001101001111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel89[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel89_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel89 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b10111101101111001011100111110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel89[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel89_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel89 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b10111110110100100101010111101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel89[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel89_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel89 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b10111110110101011111100111100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel89[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel89_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel89 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111110101000110110011000101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel89[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel89_Valid_Out)
	);
	Adder_64input add_k89(
		.Data1(Data_Out_Kernel89[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel89[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel89[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel89[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel89[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel89[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel89[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel89[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel89[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel89[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel89[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel89[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel89[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel89[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel89[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel89[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel89[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel89[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel89[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel89[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel89[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel89[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel89[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel89[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel89[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel89[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel89[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel89[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel89[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel89[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel89[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel89[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel89[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel89[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel89[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel89[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel89[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel89[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel89[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel89[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel89[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel89[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel89[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel89[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel89[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel89[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel89[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel89[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel89[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel89[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel89[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel89[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel89[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel89[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel89[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel89[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel89[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel89[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel89[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel89[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel89[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel89[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel89[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel89[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel89),
		.Data_Out(add_k89_Data_Out),
		.Valid_Out(add_kernel89_Valid_Out)
	);
	Batch_Norm bn_kernel89(
		.Data_A(32'b00111110000011111100010110111000),
		.Data_B(32'b00111111010111100001000010010111),
		.Data_In(add_k89_Data_Out),
		.Valid_In(add_kernel89_Valid_Out),
		.Data_Out(bn89_Data_Out),
		.Valid_Out(bn89_Valid_Out)
	);
	Relu_Core rl_kernel89(
		.Data_In(bn89_Data_Out),
		.Valid_In(bn89_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*89-1:DATA_WIDHT*88]),
		.Valid_Out(rl89_Valid_Out)
	);
//////////KERNEL90//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel90 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111111000100110111111110101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel90[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel90_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel90 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111101101000101110000111101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel90[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel90_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel90 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110001001001110100000110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel90[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel90_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel90 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111111000000001001100001001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel90[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel90_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel90 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111101000000101010110111001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel90[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel90_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel90 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110010110000101101000110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel90[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel90_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel90 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111100111010100111101010011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel90[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel90_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel90 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111101101101111001001101101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel90[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel90_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel90 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110001010011111100101100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel90[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel90_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel90 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111101110000101011011111111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel90[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel90_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel90 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110000000001001100111111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel90[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel90_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel90 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111100110001010010010011001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel90[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel90_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel90 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110010110001100011000111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel90[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel90_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel90 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111101011111010001111011001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel90[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel90_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel90 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110001011010001011111001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel90[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel90_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel90 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111100100111011111001110001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel90[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel90_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel90 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110111011000110011010000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel90[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel90_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel90 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110001000101110001111100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel90[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel90_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel90 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110001100101011100010000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel90[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel90_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel90 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110010101110101100110101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel90[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel90_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel90 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110100000001100101110100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel90[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel90_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel90 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111110001001100000010100101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel90[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel90_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel90 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111111000001101000101000001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel90[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel90_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel90 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111110001101011011001111010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel90[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel90_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel90 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111110100011001110101110001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel90[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel90_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel90 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110101001001001010011101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel90[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel90_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel90 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110001000000000010111000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel90[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel90_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel90 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111011110111010011110011110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel90[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel90_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel90 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111110100010001001011110101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel90[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel90_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel90 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111110101001001001101111100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel90[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel90_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel90 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111101100010000001101110001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel90[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel90_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel90 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110110101000011110101101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel90[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel90_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel90 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111110101000100100001010101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel90[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel90_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel90 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b00111101111000000000000000000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel90[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel90_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel90 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111110110110111001111100100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel90[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel90_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel90 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b10111110000110100101000111110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel90[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel90_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel90 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111110101111101001110100100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel90[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel90_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel90 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b00111101000010000001101001110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel90[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel90_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel90 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b00111110101100011001110110111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel90[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel90_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel90 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111110001110010100110010011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel90[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel90_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel90 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111111000111100100100001110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel90[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel90_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel90 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111110110000010001101101000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel90[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel90_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel90 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111110100111110001011110111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel90[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel90_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel90 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b00111101111010111011010100011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel90[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel90_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel90 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111111000000001101100110010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel90[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel90_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel90 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111110010100111011100011110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel90[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel90_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel90 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111101100101000101110101110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel90[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel90_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel90 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111110001110000101010111111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel90[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel90_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel90 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111110000000110100111110111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel90[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel90_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel90 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111110000001101101001000010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel90[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel90_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel90 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111110111011011010010010000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel90[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel90_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel90 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111101100100000011110111011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel90[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel90_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel90 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111101110001000110011010001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel90[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel90_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel90 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111110111011011001001111000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel90[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel90_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel90 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111110100010111111111111101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel90[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel90_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel90 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111101010100011010110111010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel90[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel90_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel90 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111110011010110011010000110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel90[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel90_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel90 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111110001001110110001111000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel90[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel90_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel90 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111110100000100100011111000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel90[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel90_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel90 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111110011011110100101001000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel90[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel90_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel90 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111110101011000011011100000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel90[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel90_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel90 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111101001111101101010001110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel90[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel90_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel90 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111110010000000110000000010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel90[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel90_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel90 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b10111101111010011000011101101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel90[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel90_Valid_Out)
	);
	Adder_64input add_k90(
		.Data1(Data_Out_Kernel90[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel90[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel90[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel90[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel90[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel90[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel90[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel90[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel90[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel90[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel90[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel90[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel90[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel90[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel90[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel90[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel90[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel90[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel90[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel90[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel90[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel90[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel90[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel90[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel90[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel90[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel90[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel90[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel90[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel90[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel90[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel90[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel90[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel90[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel90[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel90[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel90[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel90[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel90[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel90[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel90[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel90[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel90[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel90[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel90[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel90[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel90[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel90[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel90[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel90[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel90[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel90[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel90[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel90[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel90[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel90[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel90[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel90[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel90[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel90[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel90[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel90[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel90[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel90[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel90),
		.Data_Out(add_k90_Data_Out),
		.Valid_Out(add_kernel90_Valid_Out)
	);
	Batch_Norm bn_kernel90(
		.Data_A(32'b00111110001100101111010010000011),
		.Data_B(32'b10111111001110111010111111111111),
		.Data_In(add_k90_Data_Out),
		.Valid_In(add_kernel90_Valid_Out),
		.Data_Out(bn90_Data_Out),
		.Valid_Out(bn90_Valid_Out)
	);
	Relu_Core rl_kernel90(
		.Data_In(bn90_Data_Out),
		.Valid_In(bn90_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*90-1:DATA_WIDHT*89]),
		.Valid_Out(rl90_Valid_Out)
	);
//////////KERNEL91//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel91 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111111000000010000100101001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel91[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel91_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel91 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111101101001110100111001000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel91[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel91_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel91 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110010111101000010111100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel91[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel91_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel91 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110010000000101111011001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel91[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel91_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel91 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111100110101010100110010001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel91[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel91_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel91 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111101101101011110111010111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel91[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel91_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel91 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111110001001100100111010000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel91[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel91_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel91 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111101100001111010101000000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel91[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel91_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel91 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110011110110111111011000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel91[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel91_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel91 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111110010101000010111000110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel91[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel91_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel91 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111101000101111001000011100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel91[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel91_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel91 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111101110101101101101101100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel91[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel91_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel91 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110010010111110110010001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel91[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel91_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel91 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111101110101001000101001011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel91[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel91_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel91 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110000101011010110010011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel91[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel91_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel91 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111101011010100101110101011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel91[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel91_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel91 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110101111111011110101001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel91[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel91_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel91 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111110001101010100010110011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel91[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel91_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel91 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111011110110100111000111111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel91[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel91_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel91 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110100100011111100011101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel91[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel91_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel91 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110101111000100110101000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel91[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel91_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel91 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111110000100001110010111011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel91[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel91_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel91 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110010101111101110101000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel91[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel91_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel91 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111110000010011101011000001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel91[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel91_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel91 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111110100100000101111001010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel91[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel91_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel91 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110101101010100100001011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel91[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel91_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel91 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110101101010111001101000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel91[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel91_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel91 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110101100010000111010010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel91[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel91_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel91 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111101011000100011001000111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel91[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel91_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel91 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111010111000101100000001010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel91[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel91_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel91 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111110011111100000101001000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel91[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel91_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel91 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111101101110011001001101111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel91[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel91_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel91 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111110101100100001011001100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel91[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel91_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel91 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b00111110111000101010111101001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel91[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel91_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel91 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111111000100011100011101110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel91[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel91_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel91 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b10111101101001111101001011100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel91[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel91_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel91 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111110101010011101001011000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel91[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel91_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel91 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111101111000001111100010000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel91[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel91_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel91 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b00111100010010101100000010111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel91[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel91_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel91 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111100011010101111010000111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel91[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel91_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel91 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111110110100100000111101111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel91[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel91_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel91 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111110011001001010011110110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel91[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel91_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel91 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b00111100000011110111011110110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel91[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel91_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel91 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111100111010111010101101011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel91[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel91_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel91 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111110100000001101010011101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel91[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel91_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel91 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111110101111010010110010100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel91[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel91_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel91 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111110101111001101111001011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel91[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel91_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel91 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111111000001111111100011100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel91[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel91_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel91 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111101010000010001100110100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel91[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel91_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel91 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b00111100111011101010100110111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel91[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel91_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel91 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b10111101101011100000001010001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel91[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel91_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel91 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111110101001111101011001001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel91[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel91_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel91 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b00111110010110001100100000101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel91[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel91_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel91 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111111000001101001000110111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel91[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel91_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel91 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111100100010110000111000101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel91[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel91_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel91 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111110100010111000010010011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel91[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel91_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel91 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111110101011000110000001000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel91[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel91_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel91 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111100100010111100101111010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel91[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel91_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel91 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b10111110010011000110010011110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel91[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel91_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel91 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b00111110000101010011010110001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel91[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel91_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel91 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111100000001101011001000010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel91[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel91_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel91 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b10111101000011010110011011100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel91[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel91_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel91 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b10111100100010100111101011001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel91[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel91_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel91 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b10111101101001001110111010001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel91[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel91_Valid_Out)
	);
	Adder_64input add_k91(
		.Data1(Data_Out_Kernel91[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel91[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel91[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel91[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel91[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel91[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel91[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel91[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel91[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel91[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel91[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel91[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel91[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel91[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel91[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel91[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel91[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel91[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel91[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel91[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel91[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel91[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel91[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel91[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel91[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel91[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel91[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel91[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel91[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel91[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel91[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel91[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel91[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel91[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel91[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel91[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel91[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel91[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel91[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel91[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel91[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel91[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel91[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel91[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel91[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel91[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel91[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel91[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel91[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel91[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel91[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel91[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel91[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel91[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel91[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel91[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel91[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel91[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel91[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel91[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel91[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel91[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel91[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel91[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel91),
		.Data_Out(add_k91_Data_Out),
		.Valid_Out(add_kernel91_Valid_Out)
	);
	Batch_Norm bn_kernel91(
		.Data_A(32'b00111110010010111111101110101100),
		.Data_B(32'b10111110101000111110010010011101),
		.Data_In(add_k91_Data_Out),
		.Valid_In(add_kernel91_Valid_Out),
		.Data_Out(bn91_Data_Out),
		.Valid_Out(bn91_Valid_Out)
	);
	Relu_Core rl_kernel91(
		.Data_In(bn91_Data_Out),
		.Valid_In(bn91_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*91-1:DATA_WIDHT*90]),
		.Valid_Out(rl91_Valid_Out)
	);
//////////KERNEL92//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel92 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111101111000000111001001100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel92[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel92_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel92 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110101111110101001011010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel92[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel92_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel92 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110100010110001111011011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel92[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel92_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel92 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110000011100010101111111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel92[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel92_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel92 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111110010101111110010111101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel92[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel92_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel92 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111101011101111011010100000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel92[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel92_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel92 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111111000001101110100000001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel92[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel92_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel92 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111011010101001000000111001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel92[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel92_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel92 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111111001010111100111101000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel92[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel92_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel92 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111101000000110101101111011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel92[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel92_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel92 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110010001100111010010111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel92[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel92_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel92 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111110101011101011000010001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel92[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel92_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel92 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110010001011110000010111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel92[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel92_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel92 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111110100010110111100011011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel92[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel92_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel92 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111101101110100111110001100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel92[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel92_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel92 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111110001100010100100001000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel92[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel92_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel92 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110101011101000011101110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel92[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel92_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel92 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111101100110010111101000001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel92[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel92_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel92 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111110100001100101010101000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel92[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel92_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel92 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110011000111111100101011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel92[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel92_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel92 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110111110110100011001000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel92[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel92_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel92 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111110010111001001111110001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel92[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel92_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel92 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110110101110101110001011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel92[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel92_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel92 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111111001111111110001100100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel92[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel92_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel92 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111110001101011100110101010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel92[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel92_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel92 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111101101100010101101000000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel92[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel92_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel92 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111111000001111100111000000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel92[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel92_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel92 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110011111011001111100111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel92[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel92_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel92 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111101010011010000011010100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel92[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel92_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel92 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111101110100000101100010111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel92[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel92_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel92 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111110111100110110000100110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel92[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel92_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel92 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111101111010110101001001111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel92[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel92_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel92 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111111010110000000010111110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel92[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel92_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel92 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b00111110101111111111111101010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel92[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel92_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel92 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111111000100010001010001110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel92[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel92_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel92 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b10111101001010100100101010000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel92[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel92_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel92 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111110111111111000100100010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel92[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel92_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel92 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111110101001110001001110011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel92[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel92_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel92 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b00111101111111111010101111100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel92[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel92_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel92 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111001011101100101111001010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel92[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel92_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel92 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111111000110101001001111011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel92[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel92_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel92 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111101100001011100010011010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel92[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel92_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel92 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111101010101101001111110111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel92[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel92_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel92 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b00111101101010010011011111010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel92[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel92_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel92 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111110111111111110000100101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel92[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel92_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel92 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111111001011000000010100001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel92[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel92_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel92 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111110100000111111100110000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel92[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel92_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel92 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111110101001000011101111010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel92[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel92_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel92 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111110001101010000100000111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel92[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel92_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel92 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111110000000100101111101001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel92[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel92_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel92 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111101100100111010011000100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel92[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel92_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel92 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111110110101100101010111110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel92[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel92_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel92 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111101110100010101011001001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel92[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel92_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel92 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111111001111011111010010111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel92[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel92_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel92 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111101110010011011010100001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel92[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel92_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel92 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111110111100010000011111100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel92[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel92_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel92 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111110000101011101010010100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel92[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel92_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel92 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111110000100100101111111100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel92[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel92_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel92 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b10111110010011001000111100100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel92[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel92_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel92 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b00111110011110001110101110101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel92[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel92_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel92 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111110010011111101110111000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel92[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel92_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel92 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b10111110011101100110010001000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel92[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel92_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel92 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b10111101001011001010111011001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel92[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel92_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel92 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111110100000000100111101000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel92[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel92_Valid_Out)
	);
	Adder_64input add_k92(
		.Data1(Data_Out_Kernel92[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel92[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel92[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel92[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel92[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel92[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel92[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel92[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel92[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel92[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel92[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel92[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel92[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel92[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel92[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel92[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel92[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel92[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel92[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel92[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel92[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel92[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel92[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel92[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel92[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel92[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel92[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel92[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel92[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel92[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel92[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel92[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel92[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel92[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel92[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel92[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel92[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel92[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel92[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel92[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel92[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel92[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel92[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel92[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel92[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel92[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel92[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel92[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel92[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel92[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel92[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel92[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel92[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel92[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel92[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel92[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel92[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel92[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel92[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel92[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel92[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel92[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel92[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel92[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel92),
		.Data_Out(add_k92_Data_Out),
		.Valid_Out(add_kernel92_Valid_Out)
	);
	Batch_Norm bn_kernel92(
		.Data_A(32'b00111110000001111000000010111010),
		.Data_B(32'b00111101111011011011011110110101),
		.Data_In(add_k92_Data_Out),
		.Valid_In(add_kernel92_Valid_Out),
		.Data_Out(bn92_Data_Out),
		.Valid_Out(bn92_Valid_Out)
	);
	Relu_Core rl_kernel92(
		.Data_In(bn92_Data_Out),
		.Valid_In(bn92_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*92-1:DATA_WIDHT*91]),
		.Valid_Out(rl92_Valid_Out)
	);
//////////KERNEL93//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel93 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111101100000101011010100000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel93[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel93_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel93 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111110100010000010110111000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel93[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel93_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel93 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110011111010100010101001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel93[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel93_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel93 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110100100000011101010111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel93[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel93_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel93 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111100101101000011100001001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel93[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel93_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel93 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111100000101011100011110001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel93[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel93_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel93 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111110110101101001101111101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel93[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel93_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel93 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111110100001100101110010010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel93[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel93_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel93 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111110000010011000110010111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel93[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel93_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel93 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110101010000101101010101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel93[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel93_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel93 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111101010001010100001110010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel93[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel93_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel93 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110100011011010101010001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel93[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel93_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel93 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110000000001001100011001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel93[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel93_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel93 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111110101011101110010101000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel93[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel93_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel93 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110100001100010011001001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel93[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel93_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel93 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111110011111010111010010011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel93[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel93_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel93 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111110111100001000011101100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel93[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel93_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel93 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111110101001010000001001011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel93[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel93_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel93 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111101100110100101010000010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel93[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel93_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel93 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110001000100001011100100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel93[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel93_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel93 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110101011010001011011110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel93[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel93_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel93 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111101101001110111101111000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel93[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel93_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel93 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111110110100111011010110101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel93[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel93_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel93 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111110101111110010100010001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel93[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel93_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel93 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111101000001100101111111100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel93[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel93_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel93 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111100111001010100011011111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel93[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel93_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel93 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111110100011111111000000011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel93[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel93_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel93 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111111000001111111001010011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel93[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel93_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel93 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111110000100110110101101010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel93[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel93_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel93 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110110110111001001000100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel93[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel93_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel93 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111110101000111011010011001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel93[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel93_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel93 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111110001000011011010101011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel93[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel93_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel93 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b00111110000011111101000011111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel93[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel93_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel93 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111111010010110101100011001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel93[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel93_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel93 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111110111010001110110000111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel93[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel93_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel93 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111110100111001111011111000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel93[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel93_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel93 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b10111110110110001110001001111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel93[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel93_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel93 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b00111100110111101000111101010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel93[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel93_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel93 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111110101000011001010110101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel93[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel93_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel93 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b00111110000110111100011000011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel93[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel93_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel93 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b10111111001001001000110101111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel93[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel93_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel93 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111110011001000110101000101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel93[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel93_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel93 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b00111101101011101010011111000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel93[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel93_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel93 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111011001001110010110111100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel93[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel93_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel93 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b00111110110110111010111001000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel93[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel93_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel93 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b10111110011100000010001100101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel93[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel93_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel93 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b10111110110000100110111011010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel93[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel93_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel93 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b00111110110100111111001001000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel93[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel93_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel93 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b00111101110101010101000000001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel93[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel93_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel93 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111100100100001010001010111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel93[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel93_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel93 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111101101011010111110011001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel93[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel93_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel93 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b10111110101001001100101000011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel93[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel93_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel93 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111110101010001011011001110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel93[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel93_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel93 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b00111110011110101111110111111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel93[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel93_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel93 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b10111110011110101001101010011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel93[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel93_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel93 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111010111011000001100100011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel93[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel93_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel93 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b10111110111100000000110000001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel93[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel93_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel93 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b10111110101001101000100110011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel93[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel93_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel93 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111110101100100100010000110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel93[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel93_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel93 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111110111111110111001011101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel93[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel93_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel93 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111101001111101110010110100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel93[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel93_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel93 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111110010100010101011110011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel93[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel93_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel93 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b10111110011011100001001111100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel93[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel93_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel93 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111011110100101111001000101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel93[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel93_Valid_Out)
	);
	Adder_64input add_k93(
		.Data1(Data_Out_Kernel93[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel93[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel93[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel93[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel93[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel93[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel93[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel93[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel93[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel93[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel93[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel93[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel93[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel93[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel93[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel93[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel93[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel93[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel93[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel93[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel93[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel93[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel93[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel93[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel93[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel93[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel93[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel93[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel93[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel93[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel93[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel93[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel93[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel93[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel93[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel93[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel93[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel93[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel93[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel93[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel93[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel93[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel93[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel93[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel93[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel93[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel93[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel93[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel93[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel93[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel93[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel93[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel93[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel93[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel93[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel93[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel93[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel93[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel93[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel93[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel93[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel93[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel93[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel93[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel93),
		.Data_Out(add_k93_Data_Out),
		.Valid_Out(add_kernel93_Valid_Out)
	);
	Batch_Norm bn_kernel93(
		.Data_A(32'b00111110000110100000100100100011),
		.Data_B(32'b00111110111001001011010010100001),
		.Data_In(add_k93_Data_Out),
		.Valid_In(add_kernel93_Valid_Out),
		.Data_Out(bn93_Data_Out),
		.Valid_Out(bn93_Valid_Out)
	);
	Relu_Core rl_kernel93(
		.Data_In(bn93_Data_Out),
		.Valid_In(bn93_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*93-1:DATA_WIDHT*92]),
		.Valid_Out(rl93_Valid_Out)
	);
//////////KERNEL94//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel94 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111110011011001111001000011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel94[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel94_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel94 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111101111000011001101010000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel94[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel94_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel94 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110101101001101101000101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel94[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel94_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel94 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111101000100011110011010101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel94[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel94_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel94 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111110000110011101000110101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel94[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel94_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel94 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111110111100101111000100001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel94[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel94_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel94 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111101110110101001001000110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel94[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel94_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel94 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111110010011010100111111010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel94[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel94_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel94 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111110100001111110101100011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel94[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel94_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel94 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111110011100001010110100110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel94[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel94_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel94 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111010111110001101011110001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel94[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel94_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel94 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110011000001010011010010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel94[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel94_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel94 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111110111011111110110000111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel94[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel94_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel94 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111111010010111011011101100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel94[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel94_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel94 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110111000100011111011110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel94[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel94_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel94 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111110110011111010001000001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel94[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel94_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel94 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111111001010101100010011001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel94[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel94_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel94 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111101110001100110001101010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel94[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel94_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel94 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111110110011110111011001111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel94[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel94_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel94 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110010010001110011001000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel94[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel94_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel94 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110111000011011110111110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel94[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel94_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel94 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111110001110111110101101000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel94[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel94_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel94 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111111001101000110111010001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel94[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel94_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel94 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111110100110001010100111001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel94[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel94_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel94 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111110110010010011011100101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel94[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel94_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel94 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111111000000100010101101010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel94[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel94_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel94 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111101101000011011110111111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel94[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel94_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel94 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111111000000000111111010101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel94[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel94_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel94 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111110011110111101010100101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel94[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel94_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel94 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111110000011011001000001000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel94[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel94_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel94 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111011010010000001100010100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel94[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel94_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel94 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110001111010011110001001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel94[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel94_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel94 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b00111110000110101011110000001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel94[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel94_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel94 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111110010100011110010000011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel94[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel94_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel94 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111010010110001000010010010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel94[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel94_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel94 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b10111110000000010010111001010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel94[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel94_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel94 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b10111111001011100100000111000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel94[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel94_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel94 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b00111110000010100010011001110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel94[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel94_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel94 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111110101001111000111100010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel94[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel94_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel94 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b00111101100101001111011101101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel94[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel94_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel94 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b10111111001010000010110001100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel94[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel94_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel94 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111101101011110011001000001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel94[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel94_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel94 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111110000000100100001100101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel94[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel94_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel94 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111110101110010101101101001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel94[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel94_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel94 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b00111110010110110001011111111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel94[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel94_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel94 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b10111101110010001100100000001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel94[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel94_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel94 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b10111101110100011111100010101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel94[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel94_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel94 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111110010101001111111011011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel94[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel94_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel94 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b00111110001111101111011001000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel94[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel94_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel94 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b00111110101110101101010111010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel94[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel94_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel94 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b10111111000101000111010101000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel94[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel94_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel94 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b10111101000010100000111100101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel94[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel94_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel94 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b00111110001101111111101010011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel94[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel94_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel94 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b00111110110000101111100100101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel94[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel94_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel94 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b10111110111100010101110011100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel94[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel94_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel94 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111110100100011011101110011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel94[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel94_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel94 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b10111110011011110011110101101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel94[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel94_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel94 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b10111111000001001100001001111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel94[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel94_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel94 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111110011101011011011111011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel94[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel94_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel94 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111111001000011011110110101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel94[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel94_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel94 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b10111110110100101000111011101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel94[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel94_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel94 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111101101110101010011011101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel94[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel94_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel94 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b10111111000001001110011001111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel94[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel94_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel94 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111110111010001001011010000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel94[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel94_Valid_Out)
	);
	Adder_64input add_k94(
		.Data1(Data_Out_Kernel94[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel94[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel94[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel94[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel94[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel94[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel94[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel94[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel94[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel94[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel94[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel94[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel94[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel94[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel94[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel94[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel94[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel94[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel94[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel94[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel94[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel94[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel94[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel94[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel94[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel94[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel94[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel94[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel94[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel94[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel94[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel94[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel94[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel94[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel94[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel94[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel94[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel94[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel94[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel94[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel94[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel94[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel94[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel94[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel94[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel94[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel94[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel94[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel94[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel94[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel94[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel94[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel94[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel94[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel94[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel94[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel94[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel94[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel94[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel94[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel94[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel94[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel94[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel94[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel94),
		.Data_Out(add_k94_Data_Out),
		.Valid_Out(add_kernel94_Valid_Out)
	);
	Batch_Norm bn_kernel94(
		.Data_A(32'b00111110000110101001110111010110),
		.Data_B(32'b00111110111100011000000011100000),
		.Data_In(add_k94_Data_Out),
		.Valid_In(add_kernel94_Valid_Out),
		.Data_Out(bn94_Data_Out),
		.Valid_Out(bn94_Valid_Out)
	);
	Relu_Core rl_kernel94(
		.Data_In(bn94_Data_Out),
		.Valid_In(bn94_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*94-1:DATA_WIDHT*93]),
		.Valid_Out(rl94_Valid_Out)
	);
//////////KERNEL95//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel95 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111111010010110011001010100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel95[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel95_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel95 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111110011000100001101110000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel95[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel95_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel95 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110100101011100101101000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel95[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel95_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel95 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110001111111100100000100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel95[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel95_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel95 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111101110001110100000111000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel95[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel95_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel95 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110100011100000011011100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel95[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel95_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel95 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111110000001011011011100000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel95[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel95_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel95 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111110100100010011110101110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel95[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel95_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel95 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110100001111101011010011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel95[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel95_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel95 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111110010100001101011001010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel95[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel95_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel95 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110111101101010111100011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel95[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel95_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel95 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110110111010110101110011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel95[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel95_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel95 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111110111110101100101110000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel95[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel95_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel95 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111101101001110000110111110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel95[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel95_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel95 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110010111101000010101100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel95[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel95_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel95 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111110010011010110100011101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel95[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel95_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel95 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110101011010010001101010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel95[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel95_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel95 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110000110011000110010111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel95[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel95_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel95 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110001110111011001111010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel95[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel95_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel95 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110110111101011110001011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel95[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel95_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel95 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110000011100111100110001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel95[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel95_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel95 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111111000000100011101111110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel95[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel95_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel95 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110001001001101101100100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel95[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel95_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel95 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111110111011111010011011000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel95[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel95_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel95 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111110001100001110111100010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel95[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel95_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel95 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110011001010101101110110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel95[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel95_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel95 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111101110010111110110010000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel95[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel95_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel95 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111110101100010000101000001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel95[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel95_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel95 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111100111000101010110111011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel95[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel95_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel95 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111110100010100110001000101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel95[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel95_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel95 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111110100110001100011000110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel95[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel95_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel95 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111111000010101100111100000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel95[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel95_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel95 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b00111111000111011011011011011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel95[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel95_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel95 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111101111110101111010011010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel95[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel95_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel95 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111111001100101001010110101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel95[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel95_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel95 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b10111110100001110111111111111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel95[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel95_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel95 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111100010111011001011100101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel95[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel95_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel95 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b00111110110101111001111000101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel95[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel95_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel95 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b00111110110001010110101011110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel95[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel95_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel95 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111110110000011011010111111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel95[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel95_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel95 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111111000000010010010110101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel95[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel95_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel95 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111110001110110000110000110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel95[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel95_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel95 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111110110110101000010111110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel95[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel95_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel95 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b00111110011000001101111111001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel95[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel95_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel95 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b00111110000011111111001100010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel95[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel95_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel95 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111110111011111111001100101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel95[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel95_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel95 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b10111110100001011101101001111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel95[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel95_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel95 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111110111011101000101100111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel95[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel95_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel95 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111110100110000101010011000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel95[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel95_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel95 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111110101001100010001110001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel95[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel95_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel95 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111101110110000010011001000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel95[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel95_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel95 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111110111001000011001011000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel95[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel95_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel95 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b00111100010100101111011001011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel95[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel95_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel95 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b00111101011001000001101001000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel95[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel95_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel95 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111110001011000110001111000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel95[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel95_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel95 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111110010011001101001101110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel95[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel95_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel95 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111111010001000001011110001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel95[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel95_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel95 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111110100001010110100010110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel95[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel95_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel95 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111101001100011100010000000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel95[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel95_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel95 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b00111110111100101011111101000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel95[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel95_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel95 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111100001100101001000011101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel95[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel95_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel95 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111110101101001011110000001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel95[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel95_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel95 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111110001111001011010101010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel95[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel95_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel95 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b10111110111111001011011111011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel95[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel95_Valid_Out)
	);
	Adder_64input add_k95(
		.Data1(Data_Out_Kernel95[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel95[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel95[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel95[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel95[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel95[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel95[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel95[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel95[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel95[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel95[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel95[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel95[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel95[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel95[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel95[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel95[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel95[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel95[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel95[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel95[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel95[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel95[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel95[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel95[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel95[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel95[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel95[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel95[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel95[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel95[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel95[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel95[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel95[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel95[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel95[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel95[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel95[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel95[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel95[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel95[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel95[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel95[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel95[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel95[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel95[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel95[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel95[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel95[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel95[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel95[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel95[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel95[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel95[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel95[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel95[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel95[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel95[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel95[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel95[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel95[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel95[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel95[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel95[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel95),
		.Data_Out(add_k95_Data_Out),
		.Valid_Out(add_kernel95_Valid_Out)
	);
	Batch_Norm bn_kernel95(
		.Data_A(32'b00111110001000000001101001000010),
		.Data_B(32'b10111111101001111010101100110110),
		.Data_In(add_k95_Data_Out),
		.Valid_In(add_kernel95_Valid_Out),
		.Data_Out(bn95_Data_Out),
		.Valid_Out(bn95_Valid_Out)
	);
	Relu_Core rl_kernel95(
		.Data_In(bn95_Data_Out),
		.Valid_In(bn95_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*95-1:DATA_WIDHT*94]),
		.Valid_Out(rl95_Valid_Out)
	);
//////////KERNEL96//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel96 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111111000000101100001101111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel96[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel96_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel96 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110000010001010001100101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel96[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel96_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel96 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111101100010111010101001110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel96[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel96_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel96 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110100010101111000101101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel96[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel96_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel96 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111100111100110010100111111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel96[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel96_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel96 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111101110111010000011111011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel96[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel96_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel96 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111100100000111100111111111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel96[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel96_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel96 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111110001100000101111011110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel96[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel96_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel96 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110000011101100000111000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel96[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel96_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel96 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111101001111011000111100101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel96[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel96_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel96 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111101101100000111001100001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel96[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel96_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel96 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111110011000101110100001101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel96[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel96_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel96 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111101100111101000110010000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel96[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel96_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel96 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111101100000001010000001110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel96[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel96_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel96 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110100001101101000001111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel96[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel96_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel96 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111110011011010111011011101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel96[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel96_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel96 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111111000001101101011100010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel96[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel96_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel96 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110011110110001011011000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel96[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel96_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel96 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110110101101111011001011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel96[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel96_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel96 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111100100101000100110101101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel96[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel96_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel96 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110010111011101010110000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel96[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel96_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel96 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111101100011001100101011011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel96[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel96_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel96 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110110011001111011011001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel96[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel96_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel96 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111110000011101111000001101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel96[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel96_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel96 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111100101111000011000111010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel96[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel96_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel96 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110010010011100111011011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel96[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel96_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel96 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110100001111001011001110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel96[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel96_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel96 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111110110011101100111100011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel96[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel96_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel96 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111101010100111000110001001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel96[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel96_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel96 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111110111011001111111000011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel96[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel96_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel96 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111101101101011001111011110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel96[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel96_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel96 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110100100001110101110000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel96[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel96_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel96 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b00111110000001101000100000001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel96[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel96_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel96 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111011101111010001010001100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel96[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel96_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel96 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111110101111101001101001110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel96[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel96_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel96 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b10111101010111101101100111110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel96[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel96_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel96 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111110100001111010101001001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel96[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel96_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel96 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111101010001001100010111010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel96[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel96_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel96 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b00111110100101111100111011111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel96[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel96_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel96 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111110010111011111001011011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel96[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel96_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel96 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111111001101001011110110111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel96[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel96_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel96 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111110001100011100010000110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel96[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel96_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel96 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111101100001101000001100010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel96[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel96_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel96 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111110001110011001010110101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel96[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel96_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel96 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111101110111010110111011000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel96[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel96_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel96 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111110000100111011011100101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel96[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel96_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel96 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111110101000000111101100111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel96[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel96_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel96 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111101011111000000110001111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel96[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel96_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel96 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111101010100110001101000101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel96[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel96_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel96 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111101011100001010000101001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel96[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel96_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel96 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111110101000111001011011101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel96[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel96_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel96 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b10111011110000001001011111110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel96[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel96_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel96 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111110000111101100010100100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel96[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel96_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel96 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111110100100110000111011000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel96[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel96_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel96 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111110011100101000110010111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel96[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel96_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel96 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b00111101101101010000100110011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel96[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel96_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel96 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111110011100110011110100101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel96[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel96_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel96 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111110010111000111101000001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel96[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel96_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel96 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111101101000011010100001011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel96[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel96_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel96 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111101111011000011000010000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel96[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel96_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel96 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111110001000100011100101101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel96[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel96_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel96 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111101111011101001000101000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel96[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel96_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel96 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111110101011010011111000010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel96[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel96_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel96 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b10111101101010101011010111110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel96[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel96_Valid_Out)
	);
	Adder_64input add_k96(
		.Data1(Data_Out_Kernel96[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel96[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel96[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel96[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel96[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel96[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel96[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel96[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel96[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel96[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel96[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel96[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel96[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel96[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel96[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel96[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel96[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel96[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel96[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel96[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel96[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel96[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel96[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel96[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel96[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel96[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel96[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel96[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel96[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel96[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel96[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel96[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel96[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel96[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel96[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel96[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel96[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel96[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel96[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel96[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel96[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel96[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel96[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel96[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel96[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel96[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel96[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel96[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel96[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel96[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel96[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel96[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel96[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel96[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel96[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel96[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel96[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel96[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel96[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel96[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel96[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel96[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel96[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel96[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel96),
		.Data_Out(add_k96_Data_Out),
		.Valid_Out(add_kernel96_Valid_Out)
	);
	Batch_Norm bn_kernel96(
		.Data_A(32'b00111110010111010010001001011010),
		.Data_B(32'b10111111000110010000101001011100),
		.Data_In(add_k96_Data_Out),
		.Valid_In(add_kernel96_Valid_Out),
		.Data_Out(bn96_Data_Out),
		.Valid_Out(bn96_Valid_Out)
	);
	Relu_Core rl_kernel96(
		.Data_In(bn96_Data_Out),
		.Valid_In(bn96_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*96-1:DATA_WIDHT*95]),
		.Valid_Out(rl96_Valid_Out)
	);
//////////KERNEL97//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel97 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110110011111000001011110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel97[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel97_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel97 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111101110110111111011101010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel97[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel97_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel97 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111101110001000001010011001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel97[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel97_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel97 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110110011101100110001111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel97[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel97_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel97 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111101100000101110111011100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel97[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel97_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel97 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111101001011001101100110110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel97[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel97_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel97 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111110100011011101111110101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel97[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel97_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel97 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111110001011001010011111010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel97[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel97_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel97 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111110111101010101111110110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel97[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel97_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel97 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111011011100011010111101101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel97[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel97_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel97 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110000010001111001011001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel97[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel97_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel97 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110001011111111000011101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel97[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel97_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel97 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111100000000111000011010110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel97[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel97_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel97 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111110100000111110010000100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel97[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel97_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel97 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110110001111100101000100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel97[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel97_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel97 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111101100010101001101110100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel97[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel97_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel97 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111110101011001010000110111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel97[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel97_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel97 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111101001001101011000111010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel97[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel97_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel97 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111110000101000000101001001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel97[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel97_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel97 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111110001010011110101101101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel97[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel97_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel97 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110110010000011101011001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel97[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel97_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel97 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111101101100010100110100000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel97[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel97_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel97 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111110110000001001011011010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel97[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel97_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel97 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111110011101011001100101001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel97[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel97_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel97 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111110010100100001110001001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel97[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel97_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel97 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111101111011110101000111011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel97[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel97_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel97 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111110010111100111101011100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel97[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel97_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel97 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111110110000101001110001010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel97[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel97_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel97 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111110011000000110000010001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel97[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel97_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel97 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110110001011101110000001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel97[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel97_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel97 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111100001001000000001110000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel97[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel97_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel97 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111101001100000001110101001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel97[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel97_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel97 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b00111110011101111111010000100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel97[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel97_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel97 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111110011111101000111111100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel97[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel97_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel97 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111110111111100111100011100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel97[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel97_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel97 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111110000011001010100111101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel97[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel97_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel97 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b10111110000101101010000110001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel97[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel97_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel97 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111101001100101001000011011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel97[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel97_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel97 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111110110010101100110001001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel97[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel97_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel97 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111101011001010010000110110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel97[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel97_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel97 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b10111110100010101011000111010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel97[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel97_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel97 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b10111100000100011000111000101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel97[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel97_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel97 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b00111110001111010011110010100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel97[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel97_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel97 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b00111100011110100011111111001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel97[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel97_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel97 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b00111110010111101001000010101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel97[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel97_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel97 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b10111101100011001100001111110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel97[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel97_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel97 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b10111110100100110100001111001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel97[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel97_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel97 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b00111110110101101101111011111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel97[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel97_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel97 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111101000101110101010110001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel97[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel97_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel97 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b00111101110111110101100101001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel97[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel97_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel97 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111101010111000110010000000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel97[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel97_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel97 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b10111110100011010001111101110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel97[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel97_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel97 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b00111101000110001010100111111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel97[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel97_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel97 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b00111110010001111110100101011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel97[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel97_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel97 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111101100101100111011111101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel97[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel97_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel97 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b00111101101001001011011011100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel97[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel97_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel97 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b10111110101111000001001111110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel97[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel97_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel97 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b10111110110111101111101010110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel97[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel97_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel97 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111110010010101010000001100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel97[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel97_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel97 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111100011011010101010000100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel97[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel97_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel97 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b10111110000010010011111000110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel97[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel97_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel97 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111110000010000100110001001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel97[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel97_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel97 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111101111000011110010100101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel97[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel97_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel97 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111101101010100100111100101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel97[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel97_Valid_Out)
	);
	Adder_64input add_k97(
		.Data1(Data_Out_Kernel97[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel97[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel97[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel97[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel97[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel97[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel97[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel97[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel97[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel97[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel97[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel97[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel97[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel97[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel97[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel97[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel97[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel97[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel97[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel97[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel97[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel97[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel97[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel97[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel97[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel97[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel97[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel97[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel97[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel97[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel97[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel97[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel97[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel97[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel97[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel97[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel97[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel97[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel97[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel97[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel97[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel97[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel97[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel97[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel97[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel97[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel97[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel97[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel97[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel97[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel97[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel97[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel97[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel97[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel97[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel97[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel97[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel97[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel97[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel97[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel97[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel97[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel97[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel97[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel97),
		.Data_Out(add_k97_Data_Out),
		.Valid_Out(add_kernel97_Valid_Out)
	);
	Batch_Norm bn_kernel97(
		.Data_A(32'b00111110010101101010000010010010),
		.Data_B(32'b10111100110110011010011010110101),
		.Data_In(add_k97_Data_Out),
		.Valid_In(add_kernel97_Valid_Out),
		.Data_Out(bn97_Data_Out),
		.Valid_Out(bn97_Valid_Out)
	);
	Relu_Core rl_kernel97(
		.Data_In(bn97_Data_Out),
		.Valid_In(bn97_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*97-1:DATA_WIDHT*96]),
		.Valid_Out(rl97_Valid_Out)
	);
//////////KERNEL98//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel98 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111111001110000000111110111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel98[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel98_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel98 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111110110011111011001011010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel98[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel98_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel98 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110100110001000011100111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel98[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel98_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel98 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111101111100100110011100100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel98[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel98_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel98 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111101111111101100010010000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel98[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel98_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel98 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110101001101111110010010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel98[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel98_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel98 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111110110101100100111000101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel98[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel98_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel98 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111111001010100000111010100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel98[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel98_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel98 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111101100011010011011111100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel98[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel98_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel98 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111110000011110000000001011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel98[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel98_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel98 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111110010000111010001000010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel98[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel98_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel98 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111110011000101110110010100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel98[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel98_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel98 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111111000110111110010101011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel98[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel98_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel98 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111100101101100010011010110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel98[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel98_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel98 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110101111000101100100010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel98[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel98_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel98 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111110101100011111111101110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel98[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel98_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel98 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110000011010011000110011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel98[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel98_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel98 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111101000110101111011110100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel98[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel98_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel98 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111101101001010110000110110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel98[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel98_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel98 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111101110110100111000001111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel98[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel98_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel98 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110101001010110001000101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel98[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel98_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel98 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111111010000101001100110010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel98[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel98_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel98 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110001100010101101101101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel98[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel98_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel98 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111110101101000011100010000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel98[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel98_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel98 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111111000010100011010111110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel98[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel98_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel98 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111110011001110110000110100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel98[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel98_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel98 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111101101011110100010011111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel98[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel98_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel98 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111110010000111001011110101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel98[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel98_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel98 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111110000101001111100111101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel98[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel98_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel98 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111111000101010111110001001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel98[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel98_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel98 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111110100101111110011111101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel98[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel98_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel98 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110000101110000100110010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel98[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel98_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel98 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b00111110101010010110100000001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel98[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel98_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel98 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111110100011111000001010010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel98[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel98_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel98 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111111001100010111101100110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel98[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel98_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel98 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b10111110110000000011110011100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel98[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel98_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel98 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111011010001110001111101110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel98[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel98_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel98 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b00111111001001101010100111110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel98[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel98_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel98 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b00111110110000110010111111010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel98[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel98_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel98 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111110101011110000101110010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel98[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel98_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel98 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111101001011000110010010001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel98[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel98_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel98 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b10111101110111111010101000111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel98[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel98_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel98 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111110000011010000111111011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel98[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel98_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel98 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b00111110100000011111101100010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel98[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel98_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel98 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b00111100100011000001100111001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel98[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel98_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel98 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111111000100101010110011000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel98[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel98_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel98 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111101100001100101010100100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel98[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel98_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel98 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111110100000000101011101001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel98[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel98_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel98 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111110111110100011110111001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel98[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel98_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel98 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111110010101101100001110001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel98[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel98_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel98 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111110010011001010000111101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel98[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel98_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel98 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111110010000100101110011101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel98[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel98_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel98 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b00111110101110101011010000010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel98[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel98_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel98 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b00111110010001001110110111010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel98[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel98_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel98 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b10111101101000011111110101011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel98[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel98_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel98 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111110110001011101000111001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel98[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel98_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel98 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111111100010110110101011001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel98[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel98_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel98 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111101101110010101010101110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel98[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel98_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel98 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111101011011110111001100101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel98[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel98_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel98 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b00111110111001011010111010010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel98[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel98_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel98 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111101110011000001100111111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel98[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel98_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel98 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111101011011010000101001110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel98[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel98_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel98 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b10111101000011001000001010001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel98[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel98_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel98 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111010011011011101111110110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel98[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel98_Valid_Out)
	);
	Adder_64input add_k98(
		.Data1(Data_Out_Kernel98[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel98[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel98[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel98[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel98[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel98[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel98[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel98[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel98[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel98[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel98[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel98[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel98[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel98[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel98[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel98[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel98[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel98[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel98[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel98[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel98[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel98[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel98[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel98[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel98[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel98[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel98[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel98[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel98[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel98[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel98[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel98[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel98[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel98[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel98[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel98[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel98[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel98[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel98[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel98[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel98[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel98[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel98[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel98[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel98[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel98[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel98[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel98[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel98[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel98[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel98[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel98[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel98[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel98[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel98[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel98[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel98[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel98[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel98[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel98[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel98[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel98[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel98[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel98[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel98),
		.Data_Out(add_k98_Data_Out),
		.Valid_Out(add_kernel98_Valid_Out)
	);
	Batch_Norm bn_kernel98(
		.Data_A(32'b00111110001100001100010011001000),
		.Data_B(32'b10111111011010101101011100001000),
		.Data_In(add_k98_Data_Out),
		.Valid_In(add_kernel98_Valid_Out),
		.Data_Out(bn98_Data_Out),
		.Valid_Out(bn98_Valid_Out)
	);
	Relu_Core rl_kernel98(
		.Data_In(bn98_Data_Out),
		.Valid_In(bn98_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*98-1:DATA_WIDHT*97]),
		.Valid_Out(rl98_Valid_Out)
	);
//////////KERNEL99//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel99 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110011010011011010000111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel99[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel99_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel99 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110110111011010100111011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel99[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel99_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel99 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111101110100000101100010010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel99[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel99_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel99 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110000111111100011011010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel99[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel99_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel99 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111101001101000110010110100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel99[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel99_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel99 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110100011011101101110110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel99[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel99_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel99 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111110100011000010010011110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel99[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel99_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel99 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111111010001010100000111000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel99[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel99_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel99 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111101110111111001011001100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel99[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel99_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel99 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110011010000011010000001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel99[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel99_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel99 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111100101000100010001000111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel99[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel99_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel99 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111101101001001101010001000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel99[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel99_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel99 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111111000000101111011000010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel99[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel99_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel99 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111101100000101000100001011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel99[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel99_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel99 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110001111111000001011110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel99[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel99_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel99 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111111000010101100100110111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel99[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel99_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel99 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110000101100111110011000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel99[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel99_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel99 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111101100010010010010000100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel99[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel99_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel99 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111110011001100001110011000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel99[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel99_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel99 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111110100011000010001010010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel99[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel99_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel99 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111111010010100000000100001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel99[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel99_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel99 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111110001100101101000101001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel99[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel99_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel99 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111111000100011100000001010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel99[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel99_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel99 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111101110011010110011001100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel99[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel99_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel99 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111110000100110100111111110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel99[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel99_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel99 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111111001110110000111011100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel99[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel99_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel99 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110000111101000101111111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel99[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel99_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel99 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110111101100101101101010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel99[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel99_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel99 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111110111000101011001100000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel99[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel99_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel99 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111110001010101111011111010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel99[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel99_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel99 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111110101100010001000001100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel99[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel99_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel99 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111111000001011110110011000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel99[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel99_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel99 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111110101101101111111001001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel99[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel99_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel99 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b00111110101001110010101111111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel99[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel99_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel99 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111011111100111001001100010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel99[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel99_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel99 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b10111110000110010010110010111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel99[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel99_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel99 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111111001001001011010001111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel99[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel99_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel99 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b00111101110001111100010001010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel99[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel99_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel99 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b00111110010110011101000000001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel99[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel99_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel99 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111110000001011100001010010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel99[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel99_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel99 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111110110010000101010000000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel99[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel99_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel99 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111110111001100011110110111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel99[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel99_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel99 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b00111100001110110110111010001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel99[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel99_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel99 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b00111110100101110110101100110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel99[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel99_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel99 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111111000010001101000110110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel99[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel99_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel99 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b10111110110111100001001000100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel99[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel99_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel99 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b10111101000100011101111111111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel99[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel99_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel99 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b00111110000000010100100101111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel99[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel99_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel99 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111110111010010110110011100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel99[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel99_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel99 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b00111110001100111000011011111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel99[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel99_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel99 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111110101111111110110101100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel99[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel99_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel99 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b10111110100101011111110100110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel99[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel99_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel99 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b00111100011011100010101010000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel99[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel99_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel99 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111110011110011110000000001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel99[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel99_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel99 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b10111101011101010111101001001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel99[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel99_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel99 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b00111111000100111111100010110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel99[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel99_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel99 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b10111110000010101110011011011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel99[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel99_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel99 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b10111010101011001101101100011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel99[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel99_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel99 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111101100000101011110010001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel99[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel99_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel99 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111111001001100000110011100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel99[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel99_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel99 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111110100000000111110100111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel99[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel99_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel99 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b10111110001110110010011110000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel99[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel99_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel99 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111111001000101001100100000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel99[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel99_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel99 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b10111111000010001100001111100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel99[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel99_Valid_Out)
	);
	Adder_64input add_k99(
		.Data1(Data_Out_Kernel99[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel99[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel99[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel99[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel99[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel99[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel99[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel99[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel99[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel99[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel99[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel99[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel99[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel99[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel99[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel99[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel99[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel99[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel99[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel99[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel99[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel99[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel99[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel99[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel99[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel99[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel99[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel99[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel99[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel99[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel99[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel99[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel99[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel99[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel99[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel99[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel99[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel99[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel99[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel99[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel99[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel99[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel99[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel99[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel99[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel99[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel99[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel99[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel99[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel99[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel99[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel99[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel99[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel99[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel99[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel99[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel99[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel99[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel99[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel99[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel99[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel99[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel99[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel99[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel99),
		.Data_Out(add_k99_Data_Out),
		.Valid_Out(add_kernel99_Valid_Out)
	);
	Batch_Norm bn_kernel99(
		.Data_A(32'b00111110010010101001110110101110),
		.Data_B(32'b00111111000110111101000011011001),
		.Data_In(add_k99_Data_Out),
		.Valid_In(add_kernel99_Valid_Out),
		.Data_Out(bn99_Data_Out),
		.Valid_Out(bn99_Valid_Out)
	);
	Relu_Core rl_kernel99(
		.Data_In(bn99_Data_Out),
		.Valid_In(bn99_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*99-1:DATA_WIDHT*98]),
		.Valid_Out(rl99_Valid_Out)
	);
//////////KERNEL100//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel100 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111110110100011101010110001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel100[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel100_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel100 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110010110011010100011111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel100[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel100_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel100 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111101001010100111111100010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel100[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel100_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel100 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111101000010101000100011100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel100[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel100_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel100 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111110010010011110111100100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel100[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel100_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel100 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111100111010111001110111000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel100[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel100_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel100 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111101100000010110010100001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel100[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel100_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel100 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111100101000010010111111110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel100[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel100_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel100 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111101101010110000000110010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel100[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel100_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel100 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111110010101101110111111001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel100[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel100_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel100 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111101100011110101110011100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel100[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel100_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel100 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110000101111100000010111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel100[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel100_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel100 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111110001000000001001110110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel100[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel100_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel100 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111110110000100010001010010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel100[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel100_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel100 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111101101100101001001111100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel100[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel100_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel100 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111110110000000011101110011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel100[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel100_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel100 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111110100101011111101101000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel100[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel100_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel100 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110110111100111010101100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel100[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel100_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel100 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110001111110110000100000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel100[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel100_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel100 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111101101111000110000010111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel100[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel100_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel100 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110100110101000110110000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel100[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel100_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel100 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111101110000001110101001011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel100[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel100_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel100 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110100000010010000101001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel100[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel100_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel100 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111101111111010101001010010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel100[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel100_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel100 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111110101110100111110101001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel100[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel100_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel100 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110100100000001011010100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel100[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel100_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel100 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111111001000010000011011001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel100[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel100_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel100 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111101111110000000010101100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel100[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel100_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel100 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111101010101110101000111001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel100[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel100_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel100 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111111000000011010100110100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel100[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel100_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel100 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111110111101011000101110110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel100[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel100_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel100 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110100110100001000001100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel100[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel100_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel100 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b00111101011100110000100001010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel100[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel100_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel100 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b00111110100010110011111111001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel100[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel100_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel100 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111110111110111101000011010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel100[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel100_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel100 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b10111101101000011011011100000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel100[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel100_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel100 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b10111100110010100101000001001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel100[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel100_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel100 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111110101001001001111011110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel100[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel100_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel100 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b00111101101001111000101110001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel100[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel100_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel100 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b00111100010101111001001100010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel100[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel100_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel100 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111111001100100010111101111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel100[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel100_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel100 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111101100000111001110111000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel100[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel100_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel100 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111011010010110100111000000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel100[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel100_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel100 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111110100000100100010000010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel100[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel100_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel100 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111110100000011110101010011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel100[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel100_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel100 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111110111000101110110011110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel100[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel100_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel100 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111101101011110111000001010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel100[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel100_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel100 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111101000010011010010111011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel100[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel100_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel100 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111101001011001010000000010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel100[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel100_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel100 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111110001001101010001110010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel100[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel100_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel100 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111101110001111010000110111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel100[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel100_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel100 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111110010011100011001011101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel100[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel100_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel100 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b00111110100110010101000000110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel100[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel100_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel100 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111110011111000011011111001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel100[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel100_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel100 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111110110011011100001011010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel100[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel100_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel100 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111110100010011000101010110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel100[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel100_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel100 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111110010011111100101111100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel100[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel100_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel100 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111110111010000000011000000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel100[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel100_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel100 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b10111110001111010110100010010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel100[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel100_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel100 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111100100000011111000110111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel100[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel100_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel100 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b10111101001110101010000110101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel100[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel100_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel100 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111101101011110000100001110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel100[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel100_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel100 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111111010011101000000011100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel100[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel100_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel100 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b10111110001010101111001001011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel100[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel100_Valid_Out)
	);
	Adder_64input add_k100(
		.Data1(Data_Out_Kernel100[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel100[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel100[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel100[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel100[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel100[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel100[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel100[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel100[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel100[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel100[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel100[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel100[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel100[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel100[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel100[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel100[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel100[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel100[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel100[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel100[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel100[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel100[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel100[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel100[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel100[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel100[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel100[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel100[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel100[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel100[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel100[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel100[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel100[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel100[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel100[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel100[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel100[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel100[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel100[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel100[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel100[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel100[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel100[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel100[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel100[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel100[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel100[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel100[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel100[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel100[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel100[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel100[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel100[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel100[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel100[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel100[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel100[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel100[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel100[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel100[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel100[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel100[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel100[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel100),
		.Data_Out(add_k100_Data_Out),
		.Valid_Out(add_kernel100_Valid_Out)
	);
	Batch_Norm bn_kernel100(
		.Data_A(32'b00111110011101110011100000110101),
		.Data_B(32'b10111100110000001000001110011001),
		.Data_In(add_k100_Data_Out),
		.Valid_In(add_kernel100_Valid_Out),
		.Data_Out(bn100_Data_Out),
		.Valid_Out(bn100_Valid_Out)
	);
	Relu_Core rl_kernel100(
		.Data_In(bn100_Data_Out),
		.Valid_In(bn100_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*100-1:DATA_WIDHT*99]),
		.Valid_Out(rl100_Valid_Out)
	);
//////////KERNEL101//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel101 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111101000000000100101011111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel101[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel101_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel101 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111110011001101100110000011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel101[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel101_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel101 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110010001101011011011111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel101[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel101_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel101 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110100111010000001111001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel101[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel101_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel101 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111101101110101100100000110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel101[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel101_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel101 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111101100000100001110000000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel101[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel101_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel101 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111110100001010101010001011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel101[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel101_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel101 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111110000100010011101011110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel101[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel101_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel101 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111110011001011101001111111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel101[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel101_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel101 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111101110111011110010000111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel101[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel101_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel101 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110000001110110110100010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel101[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel101_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel101 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111101101010110011000001000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel101[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel101_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel101 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111101100111010100000011010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel101[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel101_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel101 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111110011011010001111001000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel101[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel101_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel101 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110011101011100011000011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel101[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel101_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel101 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111110011110101111010011011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel101[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel101_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel101 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111110111101000000111111010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel101[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel101_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel101 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111110011100100100111100110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel101[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel101_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel101 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111101000101100010111010101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel101[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel101_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel101 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110000100011110110110011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel101[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel101_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel101 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110101010001111111000110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel101[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel101_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel101 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111100101011000000100100111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel101[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel101_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel101 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111110011001100111010110100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel101[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel101_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel101 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111110101111110011101110010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel101[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel101_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel101 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111100101000111100110000111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel101[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel101_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel101 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111101110001001000111111101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel101[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel101_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel101 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111110101011111000110000111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel101[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel101_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel101 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111110110010011100001010011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel101[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel101_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel101 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111101011111100111100011101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel101[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel101_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel101 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110101111000100010111110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel101[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel101_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel101 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111110100111101100000100100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel101[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel101_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel101 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111110000111011010010011010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel101[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel101_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel101 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b00111110010111000110000101101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel101[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel101_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel101 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111110110011101000100001010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel101[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel101_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel101 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111111000000110111110110010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel101[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel101_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel101 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111101101100001010011010010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel101[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel101_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel101 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b10111110001011010100110000110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel101[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel101_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel101 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b00111110000001100000001100100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel101[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel101_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel101 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111111000010110001100111010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel101[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel101_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel101 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b00111110100011011100011111100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel101[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel101_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel101 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b10111111001010011101110000110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel101[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel101_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel101 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111110000000110001110000111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel101[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel101_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel101 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b00111110000001101011111110111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel101[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel101_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel101 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111100111111100101000001010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel101[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel101_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel101 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b00111111000001000111010010100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel101[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel101_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel101 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b10111110100101010111100111000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel101[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel101_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel101 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b10111110000000001101001010100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel101[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel101_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel101 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b00111110110111110111000011000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel101[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel101_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel101 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b00111110010011100111100011001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel101[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel101_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel101 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b00111110001010000001000010110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel101[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel101_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel101 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111110000001111001000001111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel101[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel101_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel101 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b10111110100111010001001001101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel101[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel101_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel101 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111110110000110101101001001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel101[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel101_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel101 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b00111110010011101111101000000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel101[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel101_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel101 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b10111101100010001011011011101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel101[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel101_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel101 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b00111110000011010111000010101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel101[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel101_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel101 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b10111110101100100010010000001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel101[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel101_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel101 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b10111111000011000001001111100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel101[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel101_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel101 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111110100111010110010111000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel101[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel101_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel101 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111110100110011011001111110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel101[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel101_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel101 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111110000010110101000100110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel101[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel101_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel101 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111110011100000110111111000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel101[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel101_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel101 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b10111110100000000101101101010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel101[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel101_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel101 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111110000011110001110111111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel101[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel101_Valid_Out)
	);
	Adder_64input add_k101(
		.Data1(Data_Out_Kernel101[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel101[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel101[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel101[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel101[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel101[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel101[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel101[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel101[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel101[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel101[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel101[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel101[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel101[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel101[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel101[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel101[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel101[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel101[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel101[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel101[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel101[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel101[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel101[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel101[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel101[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel101[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel101[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel101[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel101[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel101[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel101[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel101[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel101[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel101[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel101[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel101[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel101[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel101[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel101[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel101[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel101[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel101[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel101[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel101[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel101[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel101[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel101[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel101[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel101[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel101[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel101[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel101[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel101[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel101[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel101[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel101[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel101[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel101[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel101[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel101[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel101[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel101[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel101[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel101),
		.Data_Out(add_k101_Data_Out),
		.Valid_Out(add_kernel101_Valid_Out)
	);
	Batch_Norm bn_kernel101(
		.Data_A(32'b00111110001001100111010011001111),
		.Data_B(32'b00111100111111001100011010101001),
		.Data_In(add_k101_Data_Out),
		.Valid_In(add_kernel101_Valid_Out),
		.Data_Out(bn101_Data_Out),
		.Valid_Out(bn101_Valid_Out)
	);
	Relu_Core rl_kernel101(
		.Data_In(bn101_Data_Out),
		.Valid_In(bn101_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*101-1:DATA_WIDHT*100]),
		.Valid_Out(rl101_Valid_Out)
	);
//////////KERNEL102//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel102 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111111000011011011001011000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel102[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel102_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel102 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111101100100011010101001010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel102[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel102_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel102 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110100001110000101011011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel102[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel102_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel102 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110100100101100101110001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel102[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel102_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel102 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111101110100010110000111111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel102[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel102_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel102 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111101100010100111101100110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel102[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel102_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel102 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111110001100101110101110000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel102[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel102_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel102 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111101111111110001100100011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel102[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel102_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel102 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110101000111100101111111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel102[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel102_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel102 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111100100001001111110010101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel102[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel102_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel102 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111100100110101001011111100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel102[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel102_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel102 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111110100101010110111001000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel102[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel102_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel102 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110100101100111001110110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel102[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel102_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel102 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111011000111100110100000100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel102[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel102_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel102 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110101111110011110010001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel102[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel102_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel102 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111110100001101101111110011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel102[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel102_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel102 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110110110100001010010101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel102[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel102_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel102 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111101111000010110011000000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel102[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel102_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel102 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111101100101011000010001100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel102[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel102_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel102 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110101101110001101110111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel102[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel102_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel102 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110000110001000011100100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel102[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel102_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel102 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111100111000011110111111111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel102[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel102_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel102 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110110010000111101101011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel102[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel102_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel102 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111100110011101001001100010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel102[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel102_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel102 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111110111111100000010001000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel102[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel102_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel102 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110011011101110111100011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel102[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel102_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel102 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110001111110011011010010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel102[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel102_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel102 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110010010111111011011001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel102[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel102_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel102 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111110001000110011000110111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel102[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel102_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel102 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111101100011100100101001100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel102[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel102_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel102 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111101100011011101101100001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel102[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel102_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel102 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111100001011001101100011000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel102[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel102_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel102 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111110011001110000010101100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel102[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel102_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel102 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b00111110101011001100000110101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel102[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel102_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel102 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111110111101000100101011011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel102[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel102_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel102 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b10111101101000011001010001100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel102[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel102_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel102 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111110110010000001100011010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel102[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel102_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel102 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111101001000110100101111011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel102[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel102_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel102 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111101111101111000111000111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel102[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel102_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel102 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111100110101101100110000101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel102[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel102_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel102 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111110110010110011110011010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel102[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel102_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel102 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111110011001001000110011011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel102[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel102_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel102 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111101111000100101100100001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel102[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel102_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel102 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111110000010011010000100111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel102[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel102_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel102 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111101110000110100100100110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel102[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel102_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel102 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111110010010001001100011010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel102[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel102_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel102 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111110110111000011000000111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel102[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel102_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel102 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111110110001111011100010101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel102[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel102_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel102 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111101111110010010100101000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel102[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel102_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel102 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b00111100111101000011010101100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel102[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel102_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel102 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111101100111100001100000001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel102[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel102_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel102 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111101100101101100101010011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel102[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel102_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel102 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b00111100100001111000000000001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel102[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel102_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel102 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111110100111110000101010110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel102[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel102_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel102 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111011111110101011011011110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel102[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel102_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel102 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111100111100010010100001101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel102[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel102_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel102 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111110100101001110101101111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel102[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel102_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel102 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b10111101001011111101111110101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel102[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel102_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel102 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b10111110001100100001010100101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel102[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel102_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel102 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b00111101101001011000110000110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel102[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel102_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel102 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111110000011111011001110110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel102[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel102_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel102 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111101000001011000110100101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel102[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel102_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel102 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111100100010101101010101110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel102[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel102_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel102 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b10111110000110011001011100001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel102[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel102_Valid_Out)
	);
	Adder_64input add_k102(
		.Data1(Data_Out_Kernel102[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel102[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel102[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel102[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel102[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel102[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel102[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel102[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel102[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel102[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel102[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel102[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel102[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel102[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel102[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel102[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel102[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel102[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel102[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel102[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel102[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel102[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel102[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel102[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel102[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel102[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel102[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel102[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel102[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel102[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel102[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel102[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel102[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel102[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel102[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel102[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel102[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel102[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel102[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel102[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel102[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel102[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel102[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel102[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel102[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel102[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel102[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel102[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel102[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel102[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel102[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel102[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel102[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel102[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel102[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel102[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel102[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel102[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel102[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel102[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel102[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel102[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel102[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel102[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel102),
		.Data_Out(add_k102_Data_Out),
		.Valid_Out(add_kernel102_Valid_Out)
	);
	Batch_Norm bn_kernel102(
		.Data_A(32'b00111110011100111010110100000101),
		.Data_B(32'b10111110011010001010010110000001),
		.Data_In(add_k102_Data_Out),
		.Valid_In(add_kernel102_Valid_Out),
		.Data_Out(bn102_Data_Out),
		.Valid_Out(bn102_Valid_Out)
	);
	Relu_Core rl_kernel102(
		.Data_In(bn102_Data_Out),
		.Valid_In(bn102_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*102-1:DATA_WIDHT*101]),
		.Valid_Out(rl102_Valid_Out)
	);
//////////KERNEL103//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel103 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111101101010000111010111111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel103[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel103_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel103 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111110011111000001011010011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel103[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel103_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel103 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111111001010001001001100101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel103[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel103_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel103 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111111001100011101110111010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel103[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel103_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel103 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111110000100110010001000001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel103[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel103_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel103 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111110000010110110110001100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel103[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel103_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel103 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111110111100100101001101010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel103[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel103_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel103 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111100011110001011111011101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel103[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel103_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel103 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111110011001000011010010011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel103[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel103_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel103 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111110001011011111110011110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel103[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel103_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel103 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111101110001011111011111010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel103[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel103_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel103 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111101101011010001010101000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel103[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel103_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel103 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111100101000101000000110101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel103[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel103_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel103 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111110100000001001110111011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel103[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel103_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel103 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111100001010000101101010101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel103[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel103_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel103 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111110000011010111111111100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel103[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel103_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel103 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111111000101110010010001110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel103[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel103_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel103 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110100110101000010110001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel103[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel103_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel103 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111011111110100100010111111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel103[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel103_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel103 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111101110101100100111101100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel103[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel103_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel103 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110100100110110100010000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel103[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel103_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel103 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111110011111001110110010001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel103[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel103_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel103 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111111010100011100001101110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel103[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel103_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel103 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111110110100011010001010111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel103[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel103_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel103 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111110011000111000000101011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel103[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel103_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel103 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111111000001000011111110110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel103[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel103_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel103 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111101111011011101100100111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel103[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel103_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel103 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111101111111111001011011000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel103[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel103_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel103 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111110011010111100010001110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel103[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel103_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel103 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111110010001011101011010001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel103[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel103_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel103 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111110011100001110100110111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel103[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel103_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel103 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111111011001001001110011101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel103[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel103_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel103 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111110110001100101111110101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel103[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel103_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel103 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111110110111000100001010111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel103[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel103_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel103 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111110111000101110010001001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel103[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel103_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel103 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111110001000011111000001101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel103[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel103_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel103 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b10111111011001111110001000100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel103[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel103_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel103 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111110001011010000011101111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel103[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel103_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel103 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111111001101101110110110111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel103[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel103_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel103 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b00111110011000011110011110101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel103[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel103_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel103 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b10111111010000010100010101101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel103[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel103_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel103 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b10111101100011001101010000011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel103[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel103_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel103 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b00111110100100000100101011001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel103[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel103_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel103 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b00111101000001100000100001100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel103[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel103_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel103 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b00111110110000000000111000010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel103[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel103_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel103 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b10111101011010011011100011100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel103[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel103_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel103 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111101111001001100011000011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel103[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel103_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel103 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111100111001001101100101100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel103[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel103_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel103 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b00111110001100100100110010001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel103[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel103_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel103 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111100000011101100001101101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel103[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel103_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel103 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b10111110001001101111010101001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel103[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel103_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel103 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b10111110010001010010101001001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel103[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel103_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel103 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111110100000100000011010101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel103[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel103_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel103 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111110000100000010111010100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel103[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel103_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel103 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111101110001101100101110100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel103[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel103_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel103 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b00111100001001000011010010010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel103[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel103_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel103 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b10111110010111000011110101110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel103[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel103_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel103 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b10111100100101001001111010001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel103[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel103_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel103 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111101011111111111001101110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel103[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel103_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel103 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111101101011010011101101000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel103[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel103_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel103 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b10111101111111110001110000101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel103[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel103_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel103 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111100101001100011101000101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel103[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel103_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel103 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b10111111010100001111110011000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel103[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel103_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel103 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111111000010101101111111000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel103[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel103_Valid_Out)
	);
	Adder_64input add_k103(
		.Data1(Data_Out_Kernel103[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel103[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel103[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel103[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel103[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel103[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel103[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel103[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel103[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel103[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel103[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel103[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel103[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel103[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel103[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel103[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel103[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel103[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel103[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel103[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel103[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel103[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel103[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel103[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel103[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel103[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel103[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel103[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel103[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel103[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel103[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel103[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel103[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel103[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel103[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel103[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel103[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel103[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel103[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel103[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel103[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel103[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel103[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel103[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel103[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel103[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel103[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel103[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel103[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel103[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel103[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel103[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel103[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel103[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel103[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel103[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel103[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel103[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel103[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel103[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel103[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel103[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel103[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel103[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel103),
		.Data_Out(add_k103_Data_Out),
		.Valid_Out(add_kernel103_Valid_Out)
	);
	Batch_Norm bn_kernel103(
		.Data_A(32'b00111110000000011111011111000010),
		.Data_B(32'b00111111010110100010001000110010),
		.Data_In(add_k103_Data_Out),
		.Valid_In(add_kernel103_Valid_Out),
		.Data_Out(bn103_Data_Out),
		.Valid_Out(bn103_Valid_Out)
	);
	Relu_Core rl_kernel103(
		.Data_In(bn103_Data_Out),
		.Valid_In(bn103_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*103-1:DATA_WIDHT*102]),
		.Valid_Out(rl103_Valid_Out)
	);
//////////KERNEL104//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel104 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111110111011001110010110011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel104[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel104_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel104 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110100010010001100010111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel104[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel104_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel104 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111100111111010100010101100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel104[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel104_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel104 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110111010100010100101110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel104[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel104_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel104 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111110010110011001001100010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel104[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel104_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel104 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110001000001101101000000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel104[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel104_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel104 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111101011100111101001111000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel104[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel104_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel104 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111101001100100111101000001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel104[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel104_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel104 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110000000110010000000110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel104[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel104_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel104 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110010100011101100000101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel104[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel104_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel104 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110011010000110110011101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel104[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel104_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel104 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110101010011101011100111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel104[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel104_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel104 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110011101011111000110111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel104[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel104_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel104 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111101110110001111000010010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel104[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel104_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel104 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110001111100000111111100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel104[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel104_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel104 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111101111100110111100111111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel104[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel104_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel104 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110101000001111110100111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel104[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel104_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel104 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111101000100001010000001011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel104[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel104_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel104 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111101111111110111010100101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel104[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel104_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel104 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111100111101001110111000111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel104[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel104_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel104 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110101000110111000011110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel104[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel104_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel104 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111110000001010001100111010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel104[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel104_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel104 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110111001000010000110100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel104[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel104_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel104 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111110101010000101011111111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel104[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel104_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel104 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111110100010001111000011100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel104[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel104_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel104 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110111110100111010100101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel104[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel104_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel104 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110010000011100010111010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel104[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel104_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel104 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111110010001110110010110100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel104[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel104_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel104 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111110101000010001011011101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel104[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel104_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel104 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111110101011010111010110111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel104[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel104_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel104 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111101111101100011010010010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel104[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel104_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel104 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110111100101011001000001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel104[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel104_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel104 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111110101100000010110111001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel104[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel104_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel104 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b00111101100111010011001010101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel104[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel104_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel104 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111110110000010101110110011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel104[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel104_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel104 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111110000001111000000101011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel104[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel104_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel104 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111110011010111100110100111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel104[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel104_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel104 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b00111101000011000100010000101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel104[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel104_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel104 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b00111110111111011101001111110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel104[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel104_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel104 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111110001010000000000000000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel104[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel104_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel104 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111111010001110010110110001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel104[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel104_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel104 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111111000001011010111110111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel104[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel104_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel104 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111110100110001011100101010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel104[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel104_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel104 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b00111110001000010110110010010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel104[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel104_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel104 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111111000110111000100000101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel104[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel104_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel104 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111110011110011100110011101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel104[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel104_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel104 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111110011000001111100010011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel104[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel104_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel104 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111110010100001010110111100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel104[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel104_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel104 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111100011010000000011111011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel104[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel104_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel104 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111101111010001000101011111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel104[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel104_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel104 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111110000110100110011000011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel104[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel104_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel104 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111110011010110110001010001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel104[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel104_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel104 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111110101000011001110100001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel104[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel104_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel104 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111110110001100111011001000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel104[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel104_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel104 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111101111010100001111111010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel104[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel104_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel104 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111100000101011001011001111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel104[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel104_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel104 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111110010011011111010001010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel104[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel104_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel104 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111110100101101110011101011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel104[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel104_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel104 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111110000110001111011010111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel104[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel104_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel104 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111110110010000101001100011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel104[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel104_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel104 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111110101011001000101010100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel104[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel104_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel104 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111101000100100100110001110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel104[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel104_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel104 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111111000100000000010110011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel104[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel104_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel104 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b10111110000110011110001101010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel104[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel104_Valid_Out)
	);
	Adder_64input add_k104(
		.Data1(Data_Out_Kernel104[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel104[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel104[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel104[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel104[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel104[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel104[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel104[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel104[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel104[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel104[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel104[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel104[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel104[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel104[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel104[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel104[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel104[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel104[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel104[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel104[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel104[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel104[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel104[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel104[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel104[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel104[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel104[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel104[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel104[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel104[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel104[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel104[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel104[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel104[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel104[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel104[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel104[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel104[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel104[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel104[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel104[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel104[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel104[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel104[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel104[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel104[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel104[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel104[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel104[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel104[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel104[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel104[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel104[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel104[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel104[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel104[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel104[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel104[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel104[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel104[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel104[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel104[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel104[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel104),
		.Data_Out(add_k104_Data_Out),
		.Valid_Out(add_kernel104_Valid_Out)
	);
	Batch_Norm bn_kernel104(
		.Data_A(32'b00111110001001111001100111001001),
		.Data_B(32'b10111111001100001100000110100001),
		.Data_In(add_k104_Data_Out),
		.Valid_In(add_kernel104_Valid_Out),
		.Data_Out(bn104_Data_Out),
		.Valid_Out(bn104_Valid_Out)
	);
	Relu_Core rl_kernel104(
		.Data_In(bn104_Data_Out),
		.Valid_In(bn104_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*104-1:DATA_WIDHT*103]),
		.Valid_Out(rl104_Valid_Out)
	);
//////////KERNEL105//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel105 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111110111110111110000011011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel105[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel105_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel105 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111011111000001100111000011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel105[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel105_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel105 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111101101000001111101111100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel105[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel105_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel105 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110110011001100010101000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel105[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel105_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel105 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111100001011010010001111101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel105[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel105_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel105 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111101111100001001100101101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel105[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel105_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel105 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111110000110001101111111111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel105[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel105_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel105 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111101111010101001001111000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel105[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel105_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel105 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110000100100000001101000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel105[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel105_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel105 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111101101101101100101100011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel105[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel105_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel105 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111011101011101101111111110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel105[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel105_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel105 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111110001101001010010010001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel105[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel105_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel105 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110001010111000110110011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel105[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel105_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel105 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111110011111100000100011111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel105[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel105_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel105 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111101100010110111101001011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel105[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel105_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel105 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111101111010000011110001001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel105[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel105_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel105 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110100011010001000101101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel105[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel105_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel105 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111101100100011110111111011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel105[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel105_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel105 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110000110110100010110001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel105[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel105_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel105 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111101111011010011111111100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel105[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel105_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel105 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110111001001100010001110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel105[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel105_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel105 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111110010101111001100010101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel105[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel105_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel105 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111111001101001001110110110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel105[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel105_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel105 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111111001011110001011000110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel105[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel105_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel105 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111110111100101001111101110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel105[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel105_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel105 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110101010011000110101111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel105[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel105_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel105 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110011000110000110100011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel105[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel105_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel105 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111101111111111100111011110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel105[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel105_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel105 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111110110010010110110110111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel105[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel105_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel105 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111110101011011110110000100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel105[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel105_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel105 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111110011000110100000001010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel105[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel105_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel105 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110001110110010011101001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel105[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel105_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel105 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111111001011111001011000011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel105[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel105_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel105 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111101101111011000000110000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel105[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel105_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel105 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111110101010101101010100111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel105[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel105_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel105 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111101100001010100110101010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel105[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel105_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel105 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111110100100101111111011100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel105[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel105_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel105 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111011101100101010001110101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel105[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel105_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel105 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b00111111000010011100010010011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel105[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel105_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel105 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111110101100111010000111110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel105[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel105_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel105 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111111010100001101101000001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel105[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel105_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel105 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111110100000111011110110100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel105[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel105_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel105 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111110100101111111110011001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel105[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel105_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel105 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b00111110111000010101110010011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel105[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel105_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel105 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111111001000100011000100110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel105[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel105_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel105 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111110100100001111110101011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel105[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel105_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel105 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b10111101011000010001101010010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel105[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel105_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel105 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111101110000001111101000100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel105[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel105_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel105 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111110100100000010110100100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel105[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel105_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel105 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111110000101011000101010100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel105[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel105_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel105 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111111000001101101001101110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel105[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel105_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel105 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111110011001101000110111010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel105[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel105_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel105 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111100111101001101111100110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel105[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel105_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel105 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111111001100100100010001011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel105[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel105_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel105 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111110011110001000101010011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel105[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel105_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel105 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111101001100001110111001101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel105[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel105_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel105 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111110011111011100100011010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel105[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel105_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel105 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111110111011001111101001100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel105[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel105_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel105 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111101010011010001101000001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel105[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel105_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel105 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111110010010001110100001010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel105[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel105_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel105 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111110110110010110100101110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel105[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel105_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel105 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b10111110000100111101100111011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel105[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel105_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel105 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111111000010011011110000010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel105[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel105_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel105 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b10111100101000100101111010001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel105[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel105_Valid_Out)
	);
	Adder_64input add_k105(
		.Data1(Data_Out_Kernel105[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel105[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel105[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel105[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel105[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel105[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel105[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel105[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel105[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel105[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel105[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel105[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel105[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel105[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel105[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel105[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel105[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel105[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel105[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel105[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel105[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel105[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel105[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel105[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel105[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel105[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel105[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel105[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel105[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel105[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel105[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel105[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel105[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel105[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel105[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel105[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel105[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel105[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel105[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel105[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel105[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel105[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel105[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel105[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel105[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel105[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel105[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel105[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel105[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel105[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel105[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel105[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel105[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel105[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel105[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel105[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel105[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel105[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel105[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel105[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel105[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel105[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel105[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel105[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel105),
		.Data_Out(add_k105_Data_Out),
		.Valid_Out(add_kernel105_Valid_Out)
	);
	Batch_Norm bn_kernel105(
		.Data_A(32'b00111110000000010011010010101011),
		.Data_B(32'b10111110101000000100001010101111),
		.Data_In(add_k105_Data_Out),
		.Valid_In(add_kernel105_Valid_Out),
		.Data_Out(bn105_Data_Out),
		.Valid_Out(bn105_Valid_Out)
	);
	Relu_Core rl_kernel105(
		.Data_In(bn105_Data_Out),
		.Valid_In(bn105_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*105-1:DATA_WIDHT*104]),
		.Valid_Out(rl105_Valid_Out)
	);
//////////KERNEL106//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel106 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111101100110011001000001011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel106[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel106_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel106 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111110110100011011110111001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel106[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel106_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel106 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110010100010111111111010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel106[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel106_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel106 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110101111010010100000000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel106[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel106_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel106 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111101110011010111101101001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel106[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel106_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel106 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111101100111001011101000101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel106[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel106_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel106 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111101011011011000100111010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel106[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel106_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel106 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111101110110101100100101011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel106[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel106_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel106 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111110100010010101011010101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel106[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel106_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel106 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110010001100000000010011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel106[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel106_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel106 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110001111011110011010101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel106[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel106_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel106 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111101111111011001100001101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel106[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel106_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel106 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111101100010111011000011000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel106[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel106_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel106 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111110100011000010000010000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel106[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel106_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel106 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110010111001011010100100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel106[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel106_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel106 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111101010110110111101110000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel106[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel106_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel106 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111110001000100100111010010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel106[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel106_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel106 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111101100110100100111001011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel106[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel106_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel106 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110001100010010100001001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel106[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel106_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel106 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111101011000101101100010001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel106[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel106_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel106 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111111000001010011100010010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel106[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel106_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel106 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111110100000000001011101100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel106[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel106_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel106 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111110011100111001110101000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel106[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel106_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel106 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111110100111011000001111111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel106[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel106_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel106 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111011010001111100110000001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel106[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel106_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel106 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111101100100011100011011010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel106[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel106_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel106 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111110100010101010000011010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel106[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel106_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel106 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111111000010100110100011111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel106[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel106_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel106 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111101001111011011110101111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel106[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel106_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel106 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110100000110100110110011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel106[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel106_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel106 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111101100011110100100101010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel106[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel106_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel106 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111101101011100100000111001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel106[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel106_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel106 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b00111110101101011011110011100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel106[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel106_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel106 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111110101110111111101010011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel106[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel106_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel106 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111110111111010100010010011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel106[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel106_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel106 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111101100001111001111001101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel106[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel106_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel106 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b10111101110000000100001110110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel106[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel106_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel106 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111101110101011010101100111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel106[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel106_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel106 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111110111111101101101000100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel106[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel106_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel106 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b00111101101001111101010001111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel106[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel106_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel106 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b10111110110110011101100100110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel106[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel106_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel106 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111101101010101001010110001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel106[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel106_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel106 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111101011111010010100001111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel106[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel106_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel106 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111101111010101100001110101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel106[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel106_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel106 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b00111110101100001100011110000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel106[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel106_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel106 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b10111110110110010110011011100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel106[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel106_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel106 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111110000100101100101100001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel106[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel106_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel106 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b00111110111110100101101101100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel106[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel106_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel106 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b00111100101000100001100100010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel106[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel106_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel106 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b00111110010110011001000101011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel106[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel106_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel106 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111110101110011010000001010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel106[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel106_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel106 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b10111110100010111101010101100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel106[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel106_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel106 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111110100100100111101001001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel106[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel106_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel106 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b00111110000010110010100000110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel106[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel106_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel106 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111101100011101111111010010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel106[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel106_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel106 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b00111101111110010011100001001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel106[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel106_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel106 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b10111110110001001111000110000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel106[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel106_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel106 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b10111110111111101100110001100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel106[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel106_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel106 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111110100110000001110111000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel106[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel106_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel106 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111110100010110011100101101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel106[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel106_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel106 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111101011000110000000001011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel106[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel106_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel106 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111101111010010001111110100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel106[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel106_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel106 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b10111011101000011100001000001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel106[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel106_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel106 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111110010011000001011101011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel106[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel106_Valid_Out)
	);
	Adder_64input add_k106(
		.Data1(Data_Out_Kernel106[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel106[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel106[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel106[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel106[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel106[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel106[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel106[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel106[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel106[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel106[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel106[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel106[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel106[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel106[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel106[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel106[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel106[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel106[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel106[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel106[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel106[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel106[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel106[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel106[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel106[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel106[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel106[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel106[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel106[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel106[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel106[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel106[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel106[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel106[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel106[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel106[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel106[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel106[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel106[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel106[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel106[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel106[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel106[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel106[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel106[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel106[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel106[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel106[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel106[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel106[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel106[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel106[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel106[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel106[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel106[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel106[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel106[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel106[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel106[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel106[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel106[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel106[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel106[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel106),
		.Data_Out(add_k106_Data_Out),
		.Valid_Out(add_kernel106_Valid_Out)
	);
	Batch_Norm bn_kernel106(
		.Data_A(32'b00111110010000001011111100000101),
		.Data_B(32'b00111110101101011100101110011110),
		.Data_In(add_k106_Data_Out),
		.Valid_In(add_kernel106_Valid_Out),
		.Data_Out(bn106_Data_Out),
		.Valid_Out(bn106_Valid_Out)
	);
	Relu_Core rl_kernel106(
		.Data_In(bn106_Data_Out),
		.Valid_In(bn106_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*106-1:DATA_WIDHT*105]),
		.Valid_Out(rl106_Valid_Out)
	);
//////////KERNEL107//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel107 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111101101011001011111000010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel107[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel107_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel107 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111110110100010110001000001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel107[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel107_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel107 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110010010010101010100011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel107[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel107_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel107 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111111000010001100111101001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel107[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel107_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel107 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111101100000001011001111001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel107[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel107_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel107 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111100000111101011001100101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel107[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel107_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel107 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111110010010100100100101010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel107[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel107_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel107 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111101111000011110110101111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel107[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel107_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel107 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111110100111001001010111010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel107[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel107_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel107 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111010011101000100100111000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel107[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel107_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel107 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111100110010011010110000101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel107[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel107_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel107 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110010101010011111011110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel107[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel107_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel107 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111101010001000110101110001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel107[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel107_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel107 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111110010100010000111110010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel107[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel107_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel107 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110100010111001100100101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel107[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel107_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel107 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111101000001101011100011001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel107[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel107_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel107 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111111010111011110000100001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel107[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel107_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel107 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111100111111011011011100001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel107[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel107_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel107 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111101001000011010010111001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel107[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel107_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel107 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111100110010100010010001100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel107[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel107_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel107 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110010001011011110110111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel107[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel107_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel107 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111101110001100010100001011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel107[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel107_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel107 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111110101111100110011111010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel107[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel107_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel107 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111110011010111001001110001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel107[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel107_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel107 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111101100000101000100000111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel107[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel107_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel107 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111110100110101101011110010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel107[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel107_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel107 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111100110011010110000101100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel107[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel107_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel107 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111110100001000100101111111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel107[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel107_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel107 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111101010011001001100010111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel107[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel107_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel107 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111101101000110101101111101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel107[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel107_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel107 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111101011001101010100011001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel107[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel107_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel107 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111111000000111001001100011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel107[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel107_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel107 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b00111110001001001010011010101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel107[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel107_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel107 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111110110110101000010000101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel107[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel107_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel107 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111110000101110111000110010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel107[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel107_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel107 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111100101101010011001110000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel107[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel107_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel107 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b10111110111111110101001111101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel107[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel107_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel107 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111110000101010010000101111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel107[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel107_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel107 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111111000010000100010111100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel107[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel107_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel107 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b00111110100110010000001111101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel107[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel107_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel107 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b10111111011100100100111001110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel107[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel107_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel107 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b10111101010001111111111001100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel107[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel107_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel107 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b00111101000011100111001011111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel107[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel107_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel107 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b00111110000100111001101110000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel107[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel107_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel107 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b00111110111111100100100011100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel107[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel107_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel107 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b10111110001010000001010001100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel107[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel107_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel107 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b10111110001101110100010111110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel107[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel107_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel107 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b00111110100010000011011100100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel107[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel107_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel107 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b00111110011001111000010110011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel107[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel107_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel107 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111101111110000100111010011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel107[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel107_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel107 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b10111010110011001010111001100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel107[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel107_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel107 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b10111110011101001010011010001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel107[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel107_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel107 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111110010000110100100100011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel107[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel107_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel107 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b00111110001010100111111001110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel107[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel107_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel107 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111110100100001101000101011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel107[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel107_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel107 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111110010110101111010001011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel107[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel107_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel107 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b10111110010001000111011001000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel107[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel107_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel107 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b10111110100101110001011000111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel107[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel107_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel107 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111110001101101000010001111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel107[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel107_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel107 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111110100000000001000000110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel107[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel107_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel107 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b10111101100001000100110001101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel107[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel107_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel107 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111101111001101001001011110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel107[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel107_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel107 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b10111110100000011101101000011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel107[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel107_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel107 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111110000111111011000000101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel107[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel107_Valid_Out)
	);
	Adder_64input add_k107(
		.Data1(Data_Out_Kernel107[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel107[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel107[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel107[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel107[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel107[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel107[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel107[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel107[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel107[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel107[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel107[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel107[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel107[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel107[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel107[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel107[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel107[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel107[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel107[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel107[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel107[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel107[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel107[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel107[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel107[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel107[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel107[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel107[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel107[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel107[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel107[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel107[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel107[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel107[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel107[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel107[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel107[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel107[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel107[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel107[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel107[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel107[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel107[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel107[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel107[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel107[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel107[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel107[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel107[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel107[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel107[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel107[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel107[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel107[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel107[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel107[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel107[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel107[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel107[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel107[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel107[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel107[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel107[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel107),
		.Data_Out(add_k107_Data_Out),
		.Valid_Out(add_kernel107_Valid_Out)
	);
	Batch_Norm bn_kernel107(
		.Data_A(32'b00111110000111011100111110111010),
		.Data_B(32'b00111111000011111100111011000110),
		.Data_In(add_k107_Data_Out),
		.Valid_In(add_kernel107_Valid_Out),
		.Data_Out(bn107_Data_Out),
		.Valid_Out(bn107_Valid_Out)
	);
	Relu_Core rl_kernel107(
		.Data_In(bn107_Data_Out),
		.Valid_In(bn107_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*107-1:DATA_WIDHT*106]),
		.Valid_Out(rl107_Valid_Out)
	);
//////////KERNEL108//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel108 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110010111011000011111101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel108[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel108_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel108 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111101010101110111001100010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel108[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel108_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel108 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110100111011000011100101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel108[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel108_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel108 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111101101000010110110111101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel108[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel108_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel108 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111110100101111110110000011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel108[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel108_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel108 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111110110111101101111101101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel108[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel108_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel108 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111111011010001010001011001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel108[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel108_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel108 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111110001101100100010001000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel108[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel108_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel108 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110000111101110011111001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel108[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel108_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel108 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110010101010111011110000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel108[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel108_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel108 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110001111101111110001110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel108[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel108_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel108 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110100111111001111001101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel108[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel108_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel108 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111101100100011000000110000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel108[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel108_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel108 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111110011111101011111110100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel108[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel108_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel108 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111011101001110000011010110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel108[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel108_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel108 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111110100111110001001111110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel108[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel108_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel108 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111110101001001100000011001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel108[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel108_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel108 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110111001100000100011110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel108[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel108_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel108 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110101011100101110101110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel108[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel108_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel108 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110000110011001011101000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel108[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel108_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel108 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110110110001100100010110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel108[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel108_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel108 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111101101001011001011111011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel108[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel108_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel108 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111111000101010011101001101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel108[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel108_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel108 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111110010100111101100011110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel108[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel108_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel108 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111110111100010101010100101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel108[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel108_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel108 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111101110110010110110001000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel108[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel108_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel108 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111110001001011001000001110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel108[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel108_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel108 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111110100000110011010110101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel108[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel108_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel108 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111110100110100000000010101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel108[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel108_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel108 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110111101110010010000111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel108[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel108_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel108 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111110101011110110000110010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel108[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel108_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel108 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111110111010100000101110111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel108[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel108_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel108 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b00111101110101001110101111110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel108[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel108_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel108 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111110111011111000111000100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel108[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel108_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel108 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111111001010011000110001010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel108[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel108_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel108 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111110100010101011111011100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel108[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel108_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel108 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b10111111010110101010100111010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel108[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel108_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel108 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111110110100010011101100000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel108[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel108_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel108 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111110111110111010011011010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel108[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel108_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel108 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b00111110010111011001011101111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel108[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel108_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel108 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111101110000001001000110100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel108[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel108_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel108 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b10111100101001011110110101010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel108[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel108_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel108 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b00111100101000111001000010000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel108[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel108_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel108 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111110011011011111110111010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel108[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel108_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel108 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b00111110111110000011010000110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel108[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel108_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel108 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b10111101110001000001100011100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel108[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel108_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel108 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b10111100110010101011011101001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel108[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel108_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel108 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b00111110010010010110101000011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel108[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel108_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel108 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b00111110110101110111100011000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel108[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel108_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel108 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b00111100001010111000010101110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel108[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel108_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel108 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b10111110101000101101101100011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel108[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel108_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel108 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b10111110010110100111001101010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel108[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel108_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel108 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111111010010010110100010110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel108[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel108_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel108 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111110010001111000001111101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel108[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel108_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel108 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111110100101001010010110001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel108[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel108_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel108 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b00111110100010101010010100001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel108[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel108_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel108 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b10111111000110010000000101100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel108[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel108_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel108 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111110100010010100010010111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel108[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel108_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel108 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111110000010101111110111111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel108[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel108_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel108 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b00111101100010000111110011001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel108[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel108_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel108 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111000111010111101001011110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel108[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel108_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel108 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111110001100000000001011001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel108[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel108_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel108 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b10111110100110010010111000011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel108[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel108_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel108 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b10111101011011110110100111000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel108[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel108_Valid_Out)
	);
	Adder_64input add_k108(
		.Data1(Data_Out_Kernel108[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel108[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel108[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel108[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel108[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel108[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel108[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel108[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel108[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel108[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel108[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel108[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel108[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel108[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel108[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel108[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel108[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel108[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel108[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel108[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel108[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel108[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel108[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel108[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel108[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel108[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel108[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel108[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel108[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel108[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel108[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel108[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel108[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel108[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel108[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel108[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel108[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel108[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel108[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel108[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel108[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel108[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel108[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel108[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel108[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel108[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel108[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel108[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel108[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel108[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel108[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel108[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel108[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel108[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel108[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel108[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel108[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel108[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel108[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel108[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel108[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel108[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel108[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel108[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel108),
		.Data_Out(add_k108_Data_Out),
		.Valid_Out(add_kernel108_Valid_Out)
	);
	Batch_Norm bn_kernel108(
		.Data_A(32'b00111110000101000000110100111001),
		.Data_B(32'b00111101001101001101111011111000),
		.Data_In(add_k108_Data_Out),
		.Valid_In(add_kernel108_Valid_Out),
		.Data_Out(bn108_Data_Out),
		.Valid_Out(bn108_Valid_Out)
	);
	Relu_Core rl_kernel108(
		.Data_In(bn108_Data_Out),
		.Valid_In(bn108_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*108-1:DATA_WIDHT*107]),
		.Valid_Out(rl108_Valid_Out)
	);
//////////KERNEL109//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel109 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111110111001000001110011110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel109[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel109_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel109 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111110011110011010100011011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel109[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel109_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel109 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111101001010000101010110010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel109[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel109_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel109 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110011001011011011111110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel109[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel109_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel109 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111110100011000110000001001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel109[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel109_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel109 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111101101011111101111100100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel109[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel109_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel109 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111111000111111000000000010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel109[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel109_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel109 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111110111110100011101100111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel109[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel109_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel109 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111110000010100001101100000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel109[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel109_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel109 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111110101110001011101001101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel109[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel109_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel109 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110010101010011011110110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel109[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel109_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel109 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111100001011110110101011101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel109[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel109_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel109 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111110101110110010001001110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel109[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel109_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel109 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111110010110100100011101110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel109[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel109_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel109 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110001000110011001110100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel109[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel109_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel109 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111110001010111000010111101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel109[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel109_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel109 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110011011100110100000110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel109[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel109_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel109 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111101110111010110110000100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel109[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel109_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel109 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111110110101110111111101001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel109[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel109_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel109 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110100100001100011110110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel109[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel109_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel109 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110000110001010000100111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel109[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel109_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel109 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111111010111001000111001111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel109[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel109_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel109 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111101101100110000110010101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel109[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel109_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel109 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111110000000010110101111110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel109[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel109_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel109 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111110101001001101110000111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel109[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel109_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel109 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111101010010100010110010110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel109[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel109_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel109 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110110110000000011100001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel109[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel109_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel109 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111110010100111000100000100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel109[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel109_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel109 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111110001001111101110001101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel109[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel109_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel109 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111111100110011100111000011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel109[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel109_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel109 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111110001110001000101011110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel109[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel109_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel109 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111101101110000111101010111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel109[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel109_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel109 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b00111101100001000011111101111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel109[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel109_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel109 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111100000111011011110011101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel109[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel109_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel109 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111111001101011001000100001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel109[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel109_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel109 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b10111110010111001111101001111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel109[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel109_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel109 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111101100001000111000101011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel109[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel109_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel109 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b00111111010010111011101110111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel109[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel109_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel109 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b00111101111010001001000100001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel109[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel109_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel109 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111110101111000110100100101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel109[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel109_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel109 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b10111110001100011111111110000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel109[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel109_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel109 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111110000111110010100111110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel109[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel109_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel109 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111101010111100101001100000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel109[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel109_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel109 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b00111110100110001001010111110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel109[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel109_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel109 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111110011001001101001001011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel109[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel109_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel109 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111110100101100111000101111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel109[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel109_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel109 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111101110110111000111111111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel109[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel109_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel109 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111110110100110110111111101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel109[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel109_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel109 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111111000111101101101111101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel109[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel109_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel109 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b00111101110011101010111110010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel109[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel109_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel109 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111110000110000000100010110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel109[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel109_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel109 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111110110101010111001111000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel109[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel109_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel109 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b00111110101011101100111011010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel109[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel109_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel109 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b00111110101111001101010000001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel109[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel109_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel109 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b10111110010000010100100011110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel109[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel109_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel109 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111110000011110011111011111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel109[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel109_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel109 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111111001001010101000011111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel109[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel109_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel109 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111101000110111111111000000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel109[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel109_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel109 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111110110011011101101010110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel109[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel109_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel109 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111101100010100001110100111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel109[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel109_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel109 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b10111011010000111001100010011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel109[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel109_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel109 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b10111100111101100001000110101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel109[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel109_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel109 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b10111110011101111010110011000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel109[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel109_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel109 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111110110111010000111000111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel109[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel109_Valid_Out)
	);
	Adder_64input add_k109(
		.Data1(Data_Out_Kernel109[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel109[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel109[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel109[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel109[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel109[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel109[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel109[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel109[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel109[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel109[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel109[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel109[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel109[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel109[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel109[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel109[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel109[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel109[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel109[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel109[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel109[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel109[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel109[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel109[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel109[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel109[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel109[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel109[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel109[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel109[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel109[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel109[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel109[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel109[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel109[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel109[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel109[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel109[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel109[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel109[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel109[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel109[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel109[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel109[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel109[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel109[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel109[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel109[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel109[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel109[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel109[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel109[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel109[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel109[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel109[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel109[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel109[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel109[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel109[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel109[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel109[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel109[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel109[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel109),
		.Data_Out(add_k109_Data_Out),
		.Valid_Out(add_kernel109_Valid_Out)
	);
	Batch_Norm bn_kernel109(
		.Data_A(32'b00111110010101101110110010010001),
		.Data_B(32'b10111111010010010100001010010001),
		.Data_In(add_k109_Data_Out),
		.Valid_In(add_kernel109_Valid_Out),
		.Data_Out(bn109_Data_Out),
		.Valid_Out(bn109_Valid_Out)
	);
	Relu_Core rl_kernel109(
		.Data_In(bn109_Data_Out),
		.Valid_In(bn109_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*109-1:DATA_WIDHT*108]),
		.Valid_Out(rl109_Valid_Out)
	);
//////////KERNEL110//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel110 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110111101000100010101000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel110[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel110_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel110 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111101100010001010010111000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel110[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel110_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel110 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110001100000101111111010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel110[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel110_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel110 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111101100011110100100111110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel110[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel110_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel110 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111101111110100111101110000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel110[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel110_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel110 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111101111001100101101001010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel110[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel110_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel110 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111110100001000111111000101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel110[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel110_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel110 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111110100000010110000001101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel110[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel110_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel110 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111110111101001000000011110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel110[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel110_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel110 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110101101001010101010000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel110[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel110_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel110 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111110101010000110110001011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel110[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel110_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel110 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111110100110010001010000101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel110[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel110_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel110 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110001001101110101011111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel110[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel110_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel110 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111110111010001010001110100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel110[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel110_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel110 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110000111111011001111010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel110[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel110_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel110 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111111000000001001011111001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel110[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel110_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel110 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111111001100110011101100000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel110[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel110_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel110 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111101101100110111010000000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel110[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel110_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel110 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110001101000100000011000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel110[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel110_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel110 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111101100100100110100010011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel110[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel110_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel110 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110101101111010111000110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel110[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel110_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel110 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111110101010010001101101010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel110[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel110_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel110 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110000001111011000001011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel110[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel110_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel110 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111111010111001111101000010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel110[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel110_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel110 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111111001111110101001111111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel110[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel110_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel110 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111101010011010110010000000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel110[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel110_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel110 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111110110111101111001001100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel110[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel110_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel110 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110100100011111001010000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel110[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel110_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel110 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111101100100100000111101000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel110[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel110_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel110 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111111000010000011000100011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel110[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel110_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel110 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111100010101011011100010111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel110[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel110_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel110 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111110101111011110100001010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel110[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel110_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel110 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111100100010101000101100100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel110[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel110_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel110 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111110010111010010110111010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel110[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel110_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel110 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111111010001011000110010110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel110[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel110_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel110 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111101000111011111111011001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel110[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel110_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel110 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b10111110100001111101100101001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel110[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel110_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel110 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111111000011001110001010111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel110[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel110_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel110 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111111000010111000110010010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel110[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel110_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel110 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b00111110100101100001001110010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel110[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel110_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel110 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b10111110110110110011100001011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel110[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel110_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel110 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b10111110011110110100011100011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel110[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel110_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel110 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b00111110010001011000111111001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel110[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel110_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel110 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111110101000101001110110111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel110[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel110_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel110 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b00111110010101000110100111011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel110[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel110_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel110 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b10111111000000101001101110010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel110[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel110_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel110 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b10111100110100000011111110001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel110[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel110_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel110 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b00111111000010101011101111111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel110[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel110_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel110 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b00111110100010010000001100111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel110[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel110_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel110 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b00111101111111001011101001111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel110[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel110_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel110 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b10111011100000100110011001100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel110[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel110_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel110 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b10111110000100110010110100100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel110[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel110_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel110 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111110100000000010101111011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel110[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel110_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel110 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b00111110101100101110101100011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel110[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel110_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel110 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b10111101110010001100000101011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel110[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel110_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel110 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b00111110000111111000010101011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel110[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel110_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel110 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b10111111001111111010010011100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel110[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel110_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel110 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b10111101111100000001110010101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel110[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel110_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel110 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111101000000000011110101100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel110[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel110_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel110 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111101100001011001111111000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel110[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel110_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel110 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111101100111110110101111000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel110[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel110_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel110 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111100111010101100101110000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel110[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel110_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel110 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b10111101111011101110101100000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel110[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel110_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel110 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111110000000000110000000011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel110[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel110_Valid_Out)
	);
	Adder_64input add_k110(
		.Data1(Data_Out_Kernel110[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel110[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel110[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel110[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel110[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel110[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel110[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel110[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel110[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel110[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel110[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel110[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel110[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel110[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel110[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel110[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel110[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel110[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel110[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel110[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel110[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel110[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel110[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel110[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel110[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel110[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel110[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel110[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel110[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel110[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel110[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel110[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel110[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel110[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel110[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel110[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel110[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel110[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel110[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel110[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel110[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel110[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel110[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel110[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel110[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel110[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel110[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel110[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel110[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel110[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel110[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel110[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel110[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel110[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel110[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel110[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel110[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel110[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel110[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel110[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel110[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel110[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel110[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel110[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel110),
		.Data_Out(add_k110_Data_Out),
		.Valid_Out(add_kernel110_Valid_Out)
	);
	Batch_Norm bn_kernel110(
		.Data_A(32'b00111101111011000100011011110011),
		.Data_B(32'b00111111000111101000001011010110),
		.Data_In(add_k110_Data_Out),
		.Valid_In(add_kernel110_Valid_Out),
		.Data_Out(bn110_Data_Out),
		.Valid_Out(bn110_Valid_Out)
	);
	Relu_Core rl_kernel110(
		.Data_In(bn110_Data_Out),
		.Valid_In(bn110_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*110-1:DATA_WIDHT*109]),
		.Valid_Out(rl110_Valid_Out)
	);
//////////KERNEL111//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel111 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111110101000000101101010101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel111[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel111_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel111 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111110101011011101010111010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel111[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel111_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel111 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110000001111011011001101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel111[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel111_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel111 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110101111010011110011100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel111[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel111_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel111 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111110101110000101000001110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel111[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel111_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel111 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110001000010011111111001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel111[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel111_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel111 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111110100001100000011101011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel111[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel111_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel111 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111101101111100001100000011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel111[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel111_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel111 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111111001010111000001011000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel111[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel111_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel111 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111110100000011110100011100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel111[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel111_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel111 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111110110001101110001010101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel111[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel111_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel111 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110010000110011010101111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel111[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel111_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel111 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111110000111110111110110110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel111[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel111_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel111 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111101010110100111110110001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel111[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel111_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel111 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111101011011000001110000111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel111[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel111_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel111 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111110011000110010101100001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel111[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel111_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel111 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111110101011000010000001110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel111[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel111_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel111 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110110000111101011010111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel111[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel111_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel111 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110010010110110101011000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel111[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel111_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel111 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110101101000001000110011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel111[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel111_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel111 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111111010010001110000000110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel111[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel111_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel111 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111110010110011110100110111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel111[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel111_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel111 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111110001101000011101001101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel111[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel111_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel111 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111111010001011010101101010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel111[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel111_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel111 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111110000010011110001110011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel111[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel111_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel111 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111110100101101011011110110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel111[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel111_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel111 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111110110011111111010111010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel111[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel111_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel111 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111101001010101110001100101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel111[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel111_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel111 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111100110010110000010001001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel111[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel111_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel111 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111100101110111011101000011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel111[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel111_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel111 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111110100111010110101010011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel111[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel111_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel111 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111110100101011100110100100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel111[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel111_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel111 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b00111110110110011111011110100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel111[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel111_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel111 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111110100001101001100111001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel111[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel111_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel111 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111101111011000101101101000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel111[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel111_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel111 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b10111110000110100100010000110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel111[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel111_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel111 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b10111111001001111011100010001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel111[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel111_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel111 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b00111110011100011111101100111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel111[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel111_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel111 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111110111001000011101100110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel111[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel111_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel111 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111100011011101000001010010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel111[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel111_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel111 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b10111111011011001010000011001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel111[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel111_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel111 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b10111111000000101101010110010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel111[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel111_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel111 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b00111100101001111101101110010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel111[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel111_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel111 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111011110000010011000110111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel111[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel111_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel111 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b00111110101000110100101000101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel111[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel111_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel111 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b10111101101001011100110000000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel111[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel111_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel111 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111110100000010100010100011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel111[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel111_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel111 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b00111101110011010010001100001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel111[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel111_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel111 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111101001110010000010010110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel111[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel111_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel111 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b00111101001000100101001100111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel111[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel111_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel111 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111100000011000000100000101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel111[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel111_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel111 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111101101011010011001000001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel111[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel111_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel111 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b00111110100010010010001001101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel111[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel111_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel111 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b00111111011000010010101010011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel111[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel111_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel111 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111101100100100101111111000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel111[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel111_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel111 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b00111101101001101111101000000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel111[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel111_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel111 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111110101110101101100101010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel111[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel111_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel111 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b10111110000001001010111011100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel111[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel111_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel111 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b10111110000011111011110010011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel111[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel111_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel111 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b00111110100111000000100100011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel111[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel111_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel111 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b10111011001011100010000110100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel111[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel111_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel111 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111110101000001010001010110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel111[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel111_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel111 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b10111110110110110010110001010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel111[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel111_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel111 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111110110000010100011000001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel111[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel111_Valid_Out)
	);
	Adder_64input add_k111(
		.Data1(Data_Out_Kernel111[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel111[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel111[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel111[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel111[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel111[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel111[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel111[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel111[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel111[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel111[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel111[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel111[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel111[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel111[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel111[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel111[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel111[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel111[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel111[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel111[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel111[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel111[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel111[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel111[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel111[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel111[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel111[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel111[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel111[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel111[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel111[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel111[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel111[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel111[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel111[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel111[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel111[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel111[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel111[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel111[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel111[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel111[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel111[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel111[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel111[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel111[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel111[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel111[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel111[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel111[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel111[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel111[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel111[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel111[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel111[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel111[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel111[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel111[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel111[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel111[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel111[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel111[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel111[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel111),
		.Data_Out(add_k111_Data_Out),
		.Valid_Out(add_kernel111_Valid_Out)
	);
	Batch_Norm bn_kernel111(
		.Data_A(32'b00111110000001011001100110011101),
		.Data_B(32'b10111110001000110100111101000111),
		.Data_In(add_k111_Data_Out),
		.Valid_In(add_kernel111_Valid_Out),
		.Data_Out(bn111_Data_Out),
		.Valid_Out(bn111_Valid_Out)
	);
	Relu_Core rl_kernel111(
		.Data_In(bn111_Data_Out),
		.Valid_In(bn111_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*111-1:DATA_WIDHT*110]),
		.Valid_Out(rl111_Valid_Out)
	);
//////////KERNEL112//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel112 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111110101010010100100011011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel112[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel112_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel112 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110100000001101011100100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel112[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel112_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel112 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110101011000111010111010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel112[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel112_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel112 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110111011111001011100010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel112[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel112_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel112 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111101001100110001100000110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel112[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel112_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel112 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110000111100000001100010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel112[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel112_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel112 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111101010110011111100001100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel112[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel112_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel112 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111110000111111001111011001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel112[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel112_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel112 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111101101010110010110100101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel112[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel112_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel112 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111101100010011111100100011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel112[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel112_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel112 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110001101000000001101101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel112[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel112_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel112 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111100110100101011100000101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel112[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel112_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel112 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110001001101101101101010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel112[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel112_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel112 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111101101001000101101110100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel112[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel112_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel112 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110101011011011011011010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel112[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel112_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel112 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111110000101110110000000010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel112[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel112_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel112 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110111010101100111011011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel112[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel112_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel112 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111101110111110010011001111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel112[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel112_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel112 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111101110000101110010000000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel112[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel112_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel112 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110110001110001001000001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel112[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel112_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel112 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110110000111110101011110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel112[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel112_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel112 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111110100000011110000000101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel112[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel112_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel112 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110111010010100110110101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel112[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel112_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel112 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111110000101101111010011011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel112[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel112_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel112 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111110100001010101000010000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel112[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel112_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel112 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110100100101111000100111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel112[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel112_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel112 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110001111110011110101100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel112[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel112_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel112 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110100101000110101110100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel112[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel112_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel112 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111110101010000110111000101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel112[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel112_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel112 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111110000001010010100100111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel112[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel112_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel112 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111101000111111110010000111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel112[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel112_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel112 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110101100010010010111010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel112[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel112_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel112 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111111000001111111100101000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel112[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel112_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel112 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b00111110101011101001110010000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel112[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel112_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel112 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111110110110000101101101000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel112[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel112_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel112 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b10111110011001100111100010111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel112[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel112_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel112 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111110011001101011011011010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel112[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel112_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel112 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111101000011100000111101110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel112[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel112_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel112 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b00111101100011000101101111001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel112[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel112_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel112 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b00111100101010111111000010010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel112[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel112_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel112 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111110111101011011001100101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel112[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel112_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel112 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111110110101101011010110010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel112[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel112_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel112 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111101110001101100100000100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel112[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel112_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel112 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b00111101100011101000000001101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel112[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel112_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel112 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111110101100010110111010011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel112[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel112_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel112 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111110011000111111100001110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel112[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel112_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel112 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111110101001011001111001000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel112[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel112_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel112 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111110101100010010001000111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel112[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel112_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel112 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111110001110101111111010110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel112[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel112_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel112 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b00111110010011101010110000010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel112[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel112_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel112 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111110001110000100101011111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel112[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel112_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel112 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111110011110000001000100111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel112[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel112_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel112 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b00111101100001100110001110110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel112[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel112_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel112 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111110101101001110010111100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel112[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel112_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel112 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111100110110010111001100111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel112[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel112_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel112 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111110001010111000110110001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel112[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel112_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel112 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111110010100001001111111010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel112[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel112_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel112 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b10111101011001111010000100100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel112[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel112_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel112 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111101100101100000101110100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel112[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel112_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel112 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111100000001001111001101111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel112[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel112_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel112 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111110101110010011010100001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel112[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel112_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel112 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b10111100101001011111011101001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel112[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel112_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel112 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111101110000101010001111000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel112[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel112_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel112 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b10111101101000001111001111100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel112[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel112_Valid_Out)
	);
	Adder_64input add_k112(
		.Data1(Data_Out_Kernel112[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel112[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel112[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel112[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel112[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel112[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel112[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel112[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel112[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel112[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel112[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel112[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel112[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel112[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel112[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel112[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel112[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel112[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel112[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel112[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel112[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel112[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel112[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel112[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel112[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel112[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel112[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel112[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel112[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel112[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel112[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel112[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel112[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel112[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel112[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel112[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel112[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel112[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel112[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel112[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel112[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel112[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel112[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel112[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel112[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel112[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel112[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel112[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel112[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel112[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel112[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel112[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel112[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel112[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel112[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel112[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel112[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel112[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel112[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel112[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel112[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel112[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel112[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel112[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel112),
		.Data_Out(add_k112_Data_Out),
		.Valid_Out(add_kernel112_Valid_Out)
	);
	Batch_Norm bn_kernel112(
		.Data_A(32'b00111110010010111100111100101011),
		.Data_B(32'b10111111010101001100001111011100),
		.Data_In(add_k112_Data_Out),
		.Valid_In(add_kernel112_Valid_Out),
		.Data_Out(bn112_Data_Out),
		.Valid_Out(bn112_Valid_Out)
	);
	Relu_Core rl_kernel112(
		.Data_In(bn112_Data_Out),
		.Valid_In(bn112_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*112-1:DATA_WIDHT*111]),
		.Valid_Out(rl112_Valid_Out)
	);
//////////KERNEL113//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel113 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111110101011010110000101111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel113[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel113_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel113 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111101011111100101000001111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel113[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel113_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel113 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111101110011101000101001110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel113[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel113_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel113 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110101010101111010010100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel113[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel113_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel113 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111110000100101111000000100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel113[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel113_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel113 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110010111000100101000000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel113[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel113_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel113 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111110100010110001101010100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel113[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel113_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel113 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111101110011001100111111001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel113[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel113_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel113 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110011011000011101110111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel113[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel113_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel113 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111101110100100011000110100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel113[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel113_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel113 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111100101100001000001000110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel113[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel113_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel113 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111110000100100111011010011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel113[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel113_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel113 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110000000111101101101110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel113[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel113_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel113 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111110011001100000101011111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel113[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel113_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel113 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111101011011110111100011001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel113[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel113_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel113 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111110011010001011000001000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel113[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel113_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel113 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110010000110010101000110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel113[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel113_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel113 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111101000011000011100110010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel113[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel113_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel113 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110011010010000000110010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel113[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel113_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel113 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111110100111001100101100101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel113[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel113_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel113 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111111000000011111101110000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel113[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel113_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel113 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111110000011100111011000100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel113[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel113_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel113 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111111000010100100000001110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel113[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel113_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel113 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111110111110101000011100011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel113[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel113_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel113 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111110111011000101000100000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel113[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel113_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel113 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110111000001100001001001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel113[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel113_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel113 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110100101000111001010001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel113[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel113_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel113 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111110100100100010010110010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel113[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel113_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel113 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111111000001011011101010010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel113[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel113_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel113 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111110111100010000011111101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel113[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel113_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel113 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111100111100001111011100000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel113[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel113_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel113 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110111001011000011001011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel113[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel113_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel113 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111110110010110011110011010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel113[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel113_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel113 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111101111000101101100101001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel113[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel113_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel113 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111110000000001001110000100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel113[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel113_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel113 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111101110101010011110011111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel113[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel113_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel113 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111110101110100011001101010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel113[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel113_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel113 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b00111110011100110111001011010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel113[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel113_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel113 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b00111111001000110100011111100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel113[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel113_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel113 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111110100001011110101010111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel113[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel113_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel113 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111111010001100000011101001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel113[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel113_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel113 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111110101101010011111111001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel113[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel113_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel113 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111110100111100011010011011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel113[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel113_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel113 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b00111111001000111110000010110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel113[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel113_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel113 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111110110111000000110011101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel113[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel113_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel113 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111110010101100100110010111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel113[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel113_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel113 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b10111110100110100000110111110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel113[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel113_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel113 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111110001010010111001001010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel113[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel113_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel113 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111110110110101111110101111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel113[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel113_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel113 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111110001001011000100100001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel113[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel113_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel113 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111110101101111110011100100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel113[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel113_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel113 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111110010101110000101001011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel113[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel113_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel113 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111101011001010000001101111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel113[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel113_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel113 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111111001000110001111110010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel113[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel113_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel113 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111110000110111010111000001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel113[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel113_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel113 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b00111101000000000000111011110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel113[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel113_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel113 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111110100110100110001001010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel113[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel113_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel113 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111110110101001000000110000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel113[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel113_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel113 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111110011000101011101000011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel113[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel113_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel113 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111110110100010100101111011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel113[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel113_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel113 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111110110111000100001110111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel113[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel113_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel113 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111101001000111000111010101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel113[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel113_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel113 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111111000111011010101011000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel113[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel113_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel113 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b10111110100101100011111110111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel113[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel113_Valid_Out)
	);
	Adder_64input add_k113(
		.Data1(Data_Out_Kernel113[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel113[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel113[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel113[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel113[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel113[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel113[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel113[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel113[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel113[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel113[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel113[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel113[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel113[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel113[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel113[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel113[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel113[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel113[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel113[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel113[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel113[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel113[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel113[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel113[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel113[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel113[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel113[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel113[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel113[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel113[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel113[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel113[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel113[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel113[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel113[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel113[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel113[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel113[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel113[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel113[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel113[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel113[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel113[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel113[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel113[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel113[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel113[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel113[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel113[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel113[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel113[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel113[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel113[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel113[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel113[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel113[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel113[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel113[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel113[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel113[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel113[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel113[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel113[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel113),
		.Data_Out(add_k113_Data_Out),
		.Valid_Out(add_kernel113_Valid_Out)
	);
	Batch_Norm bn_kernel113(
		.Data_A(32'b00111110000000101011100110111000),
		.Data_B(32'b10111110011100000100100011011101),
		.Data_In(add_k113_Data_Out),
		.Valid_In(add_kernel113_Valid_Out),
		.Data_Out(bn113_Data_Out),
		.Valid_Out(bn113_Valid_Out)
	);
	Relu_Core rl_kernel113(
		.Data_In(bn113_Data_Out),
		.Valid_In(bn113_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*113-1:DATA_WIDHT*112]),
		.Valid_Out(rl113_Valid_Out)
	);
//////////KERNEL114//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel114 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111111000110011000001100001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel114[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel114_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel114 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110100000111001010110010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel114[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel114_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel114 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110100010101000100000001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel114[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel114_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel114 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110011011100011000001010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel114[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel114_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel114 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111100101011111100100011100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel114[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel114_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel114 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110001010000001110011101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel114[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel114_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel114 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111101110111110011110110110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel114[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel114_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel114 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111110100101010000110001101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel114[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel114_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel114 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110101001100101111101111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel114[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel114_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel114 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111100111000011010001010111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel114[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel114_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel114 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111101000001011010101110010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel114[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel114_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel114 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111110011010100010101111011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel114[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel114_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel114 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110000100101001110111100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel114[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel114_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel114 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111101111111110001110110110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel114[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel114_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel114 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110100101001110101101001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel114[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel114_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel114 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111101011011010110100110011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel114[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel114_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel114 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111101011001101101100111000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel114[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel114_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel114 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110100001010100001001110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel114[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel114_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel114 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110000011000011010101011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel114[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel114_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel114 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110001111001000001001101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel114[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel114_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel114 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110011110110110101010100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel114[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel114_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel114 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111100111001000110010001100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel114[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel114_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel114 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111111000100011000101010100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel114[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel114_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel114 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111101110111010011000011011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel114[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel114_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel114 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111101100000010100110000100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel114[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel114_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel114 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110100001111000010001001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel114[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel114_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel114 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110101010100010101100001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel114[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel114_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel114 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110001001010101100100010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel114[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel114_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel114 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111101111111110101111001000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel114[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel114_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel114 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111111000010011011010110100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel114[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel114_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel114 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111101101110111110110101011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel114[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel114_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel114 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111101001010111000100010010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel114[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel114_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel114 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111100100111011000101101100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel114[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel114_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel114 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b00111110011101001011011010011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel114[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel114_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel114 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111110111110100110111011101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel114[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel114_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel114 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b10111110000101100011010101000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel114[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel114_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel114 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111110100101001011100001000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel114[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel114_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel114 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111110000011000111010010101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel114[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel114_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel114 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111101111011110100010010110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel114[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel114_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel114 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111101010110110101101011011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel114[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel114_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel114 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111111000111000010011001100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel114[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel114_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel114 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111110001111011010101011100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel114[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel114_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel114 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111110001001010101010001000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel114[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel114_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel114 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111110101111001101000110111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel114[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel114_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel114 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b00111110001011000011010011010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel114[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel114_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel114 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111110001000110100100011001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel114[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel114_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel114 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111110101011101000111110111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel114[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel114_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel114 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111110000111010111011011000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel114[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel114_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel114 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111110000100100110000001011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel114[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel114_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel114 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b00111101010011110101101101001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel114[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel114_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel114 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111110001001100010100101100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel114[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel114_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel114 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b10111101100000110011001101001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel114[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel114_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel114 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111110000100110001100110011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel114[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel114_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel114 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111110001000011010010111000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel114[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel114_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel114 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111110100011011011100110001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel114[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel114_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel114 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b00111101001011100000001010010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel114[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel114_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel114 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111101000010001001001110011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel114[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel114_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel114 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111110010001001011011001001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel114[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel114_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel114 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b10111101010111111000111000010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel114[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel114_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel114 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111101000110101000111010011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel114[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel114_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel114 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111101110111101111101110101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel114[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel114_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel114 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111110000111001000011110110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel114[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel114_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel114 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111110100010101010111100011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel114[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel114_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel114 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b10111101110000110000100100010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel114[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel114_Valid_Out)
	);
	Adder_64input add_k114(
		.Data1(Data_Out_Kernel114[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel114[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel114[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel114[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel114[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel114[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel114[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel114[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel114[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel114[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel114[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel114[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel114[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel114[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel114[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel114[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel114[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel114[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel114[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel114[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel114[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel114[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel114[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel114[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel114[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel114[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel114[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel114[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel114[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel114[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel114[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel114[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel114[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel114[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel114[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel114[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel114[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel114[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel114[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel114[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel114[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel114[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel114[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel114[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel114[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel114[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel114[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel114[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel114[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel114[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel114[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel114[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel114[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel114[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel114[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel114[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel114[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel114[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel114[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel114[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel114[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel114[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel114[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel114[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel114),
		.Data_Out(add_k114_Data_Out),
		.Valid_Out(add_kernel114_Valid_Out)
	);
	Batch_Norm bn_kernel114(
		.Data_A(32'b00111110100011010010101011111011),
		.Data_B(32'b10111101111001110011111100000110),
		.Data_In(add_k114_Data_Out),
		.Valid_In(add_kernel114_Valid_Out),
		.Data_Out(bn114_Data_Out),
		.Valid_Out(bn114_Valid_Out)
	);
	Relu_Core rl_kernel114(
		.Data_In(bn114_Data_Out),
		.Valid_In(bn114_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*114-1:DATA_WIDHT*113]),
		.Valid_Out(rl114_Valid_Out)
	);
//////////KERNEL115//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel115 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110100111010100101011010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel115[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel115_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel115 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111100101010000111101101100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel115[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel115_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel115 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111101110011101010101001011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel115[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel115_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel115 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110100111001001011000000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel115[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel115_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel115 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111110001110011101010000000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel115[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel115_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel115 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111101101111101010111110010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel115[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel115_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel115 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111101010111100001111010001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel115[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel115_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel115 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111110000110111110101110000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel115[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel115_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel115 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111110101010011001110000010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel115[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel115_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel115 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111110000010010011011100100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel115[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel115_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel115 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111101001110100001010010010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel115[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel115_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel115 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111101000000001110110011110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel115[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel115_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel115 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111110000110100110111111000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel115[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel115_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel115 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111101101101010110010101000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel115[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel115_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel115 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110100011000001000000011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel115[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel115_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel115 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111110000001101011111111001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel115[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel115_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel115 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111111010101111110001100101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel115[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel115_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel115 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110011000000000000111110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel115[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel115_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel115 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111101001101001001011010001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel115[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel115_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel115 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111100110010110001101101101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel115[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel115_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel115 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111101101111101111101011001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel115[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel115_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel115 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111101010000011101111011000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel115[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel115_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel115 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111100101110011101111101001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel115[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel115_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel115 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111110011011011001000000001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel115[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel115_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel115 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111110111000110111011110110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel115[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel115_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel115 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111110100010111000001101001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel115[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel115_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel115 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111110000001001100011110000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel115[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel115_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel115 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110001101011011001010101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel115[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel115_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel115 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111101100000101100111001111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel115[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel115_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel115 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111110100010011110000110110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel115[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel115_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel115 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111110001011110101001111011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel115[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel115_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel115 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111110111000100000100010100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel115[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel115_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel115 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b00111110110110001101011101011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel115[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel115_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel115 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b00111110000000001000100010101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel115[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel115_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel115 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111110100010100001001010100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel115[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel115_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel115 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b10111101111000111101011011001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel115[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel115_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel115 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b10111111000001101010001100011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel115[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel115_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel115 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b00111101100010110001100000111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel115[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel115_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel115 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111110111100100000101100100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel115[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel115_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel115 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b00111110111010011110011100000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel115[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel115_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel115 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b10111110101001101001110110100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel115[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel115_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel115 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b10111101001101010000001011111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel115[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel115_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel115 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b00111110000000011011011011010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel115[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel115_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel115 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111101101110001110110010011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel115[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel115_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel115 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b00111110101101111010100010100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel115[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel115_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel115 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b10111101110110001100011111101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel115[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel115_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel115 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b10111110100011101100000011011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel115[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel115_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel115 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b00111110000100101011001000001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel115[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel115_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel115 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111101100101011001001000000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel115[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel115_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel115 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111110000101000000011000101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel115[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel115_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel115 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111101110011010001011001010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel115[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel115_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel115 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b10111110100100100111000000010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel115[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel115_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel115 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111110001010111011001111010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel115[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel115_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel115 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b00111110011110110011001011011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel115[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel115_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel115 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111101100011010110010001101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel115[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel115_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel115 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b00111100000011000010110010111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel115[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel115_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel115 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b10111111000000001011010011001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel115[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel115_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel115 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b10111110101110000011011111010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel115[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel115_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel115 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111101100101000001000110110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel115[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel115_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel115 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111101100010101101110010110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel115[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel115_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel115 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b10111110001100001001101100101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel115[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel115_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel115 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b10111101010110101010101001011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel115[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel115_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel115 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b10111101101000011010111100111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel115[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel115_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel115 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b10111100101110000000011100101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel115[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel115_Valid_Out)
	);
	Adder_64input add_k115(
		.Data1(Data_Out_Kernel115[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel115[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel115[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel115[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel115[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel115[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel115[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel115[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel115[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel115[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel115[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel115[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel115[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel115[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel115[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel115[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel115[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel115[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel115[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel115[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel115[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel115[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel115[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel115[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel115[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel115[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel115[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel115[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel115[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel115[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel115[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel115[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel115[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel115[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel115[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel115[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel115[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel115[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel115[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel115[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel115[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel115[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel115[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel115[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel115[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel115[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel115[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel115[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel115[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel115[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel115[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel115[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel115[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel115[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel115[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel115[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel115[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel115[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel115[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel115[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel115[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel115[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel115[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel115[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel115),
		.Data_Out(add_k115_Data_Out),
		.Valid_Out(add_kernel115_Valid_Out)
	);
	Batch_Norm bn_kernel115(
		.Data_A(32'b00111110010000101101111011011111),
		.Data_B(32'b00111110111010111111101111100011),
		.Data_In(add_k115_Data_Out),
		.Valid_In(add_kernel115_Valid_Out),
		.Data_Out(bn115_Data_Out),
		.Valid_Out(bn115_Valid_Out)
	);
	Relu_Core rl_kernel115(
		.Data_In(bn115_Data_Out),
		.Valid_In(bn115_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*115-1:DATA_WIDHT*114]),
		.Valid_Out(rl115_Valid_Out)
	);
//////////KERNEL116//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel116 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111110101110010100110001110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel116[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel116_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel116 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111101111100101001101001110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel116[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel116_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel116 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110100100111001001000011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel116[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel116_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel116 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111101110111100011000001000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel116[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel116_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel116 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111101101111000101010110001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel116[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel116_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel116 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111100000010001101010001001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel116[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel116_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel116 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111110001010111100110110010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel116[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel116_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel116 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111110001001100001010100000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel116[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel116_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel116 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111100110001000000110100101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel116[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel116_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel116 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111110011000111111111110110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel116[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel116_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel116 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111101011000010011101000100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel116[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel116_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel116 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111101110001010111111111111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel116[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel116_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel116 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111101011001101011000011001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel116[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel116_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel116 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111110001011110111110100110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel116[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel116_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel116 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111011100001001101011000101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel116[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel116_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel116 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111101110111111010111100101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel116[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel116_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel116 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110001110011111000101111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel116[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel116_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel116 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111101101001010111100110001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel116[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel116_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel116 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111101000011010010111111111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel116[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel116_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel116 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111101001000010000010111011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel116[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel116_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel116 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110001001101111010100001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel116[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel116_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel116 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111101010010100110010110001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel116[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel116_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel116 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110100010000010100100101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel116[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel116_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel116 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111101110011100011101011111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel116[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel116_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel116 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111100010000011010001101010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel116[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel116_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel116 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110010111110110100101100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel116[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel116_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel116 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110111110000100011110101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel116[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel116_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel116 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110001011101000111100100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel116[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel116_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel116 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111101110100101010100101111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel116[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel116_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel116 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111101101101011000011011011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel116[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel116_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel116 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111110101000011110110000000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel116[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel116_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel116 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110011101111000011101010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel116[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel116_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel116 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111101111110101011001000011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel116[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel116_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel116 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b00111110010000111111111100101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel116[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel116_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel116 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111110111101000101010110100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel116[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel116_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel116 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b10111101100110100110010101111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel116[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel116_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel116 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111110101011101110110111011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel116[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel116_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel116 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111110001011100011001010100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel116[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel116_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel116 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b00111110010001000101000011110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel116[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel116_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel116 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111101111000101011001101111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel116[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel116_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel116 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111111000000010010010111000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel116[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel116_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel116 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111101110110100001101110001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel116[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel116_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel116 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b00111101010101011011010101011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel116[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel116_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel116 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111101101000110000111110000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel116[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel116_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel116 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111101110110000100111011000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel116[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel116_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel116 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111110101110010110100111110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel116[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel116_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel116 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111110000011011100000100010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel116[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel116_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel116 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111110001110011000111100010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel116[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel116_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel116 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111100110111100110101100011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel116[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel116_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel116 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111101000011111111100101110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel116[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel116_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel116 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111101000111100110101111000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel116[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel116_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel116 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111110001001001011010110101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel116[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel116_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel116 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b00111110100100111111000111011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel116[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel116_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel116 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111110110011111100100011111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel116[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel116_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel116 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111110010011000010000110101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel116[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel116_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel116 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111110010011110000010101010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel116[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel116_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel116 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111110101110100101001110010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel116[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel116_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel116 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111110011100100000100001010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel116[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel116_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel116 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b10111110000001110001110010101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel116[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel116_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel116 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b00111110010111011001010000111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel116[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel116_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel116 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111101001111101101101011110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel116[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel116_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel116 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111101000010011001100010100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel116[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel116_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel116 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111110011011010011011100010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel116[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel116_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel116 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b10111101011111111000011100010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel116[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel116_Valid_Out)
	);
	Adder_64input add_k116(
		.Data1(Data_Out_Kernel116[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel116[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel116[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel116[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel116[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel116[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel116[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel116[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel116[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel116[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel116[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel116[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel116[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel116[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel116[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel116[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel116[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel116[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel116[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel116[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel116[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel116[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel116[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel116[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel116[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel116[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel116[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel116[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel116[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel116[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel116[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel116[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel116[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel116[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel116[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel116[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel116[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel116[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel116[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel116[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel116[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel116[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel116[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel116[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel116[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel116[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel116[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel116[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel116[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel116[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel116[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel116[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel116[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel116[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel116[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel116[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel116[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel116[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel116[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel116[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel116[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel116[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel116[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel116[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel116),
		.Data_Out(add_k116_Data_Out),
		.Valid_Out(add_kernel116_Valid_Out)
	);
	Batch_Norm bn_kernel116(
		.Data_A(32'b00111110011011001111100000110110),
		.Data_B(32'b10111111001111001100000011111110),
		.Data_In(add_k116_Data_Out),
		.Valid_In(add_kernel116_Valid_Out),
		.Data_Out(bn116_Data_Out),
		.Valid_Out(bn116_Valid_Out)
	);
	Relu_Core rl_kernel116(
		.Data_In(bn116_Data_Out),
		.Valid_In(bn116_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*116-1:DATA_WIDHT*115]),
		.Valid_Out(rl116_Valid_Out)
	);
//////////KERNEL117//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel117 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111101100010101101101001000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel117[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel117_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel117 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110010000111010001100001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel117[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel117_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel117 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110101110100110011010100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel117[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel117_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel117 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111111000010100011110011011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel117[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel117_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel117 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111110000001100111110100000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel117[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel117_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel117 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111101111000011111101011111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel117[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel117_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel117 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111111001111111110000001111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel117[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel117_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel117 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111101111111000000000110111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel117[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel117_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel117 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110011101011100001100111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel117[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel117_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel117 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111101100011101011000110001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel117[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel117_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel117 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111110110000000001100100011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel117[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel117_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel117 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111110110111110011011110111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel117[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel117_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel117 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110000101000110100001110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel117[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel117_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel117 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111100011011101100010011000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel117[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel117_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel117 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111101101111111000011010110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel117[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel117_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel117 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111101000000111100010100101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel117[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel117_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel117 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110111010101111111001101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel117[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel117_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel117 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111110100101111000000100110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel117[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel117_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel117 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111101101011110101011001001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel117[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel117_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel117 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111110010110010000011110001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel117[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel117_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel117 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111111000011000011011100100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel117[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel117_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel117 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111110100000111011001010110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel117[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel117_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel117 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111111010010010010111110100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel117[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel117_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel117 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111111000000010001011101011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel117[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel117_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel117 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111111000101101000010101011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel117[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel117_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel117 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111101001010001111011000110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel117[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel117_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel117 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110010111011011011101011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel117[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel117_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel117 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110000100100100111110111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel117[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel117_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel117 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111101101010001101011101001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel117[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel117_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel117 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111100001000000101011010101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel117[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel117_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel117 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111111000001011000010011110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel117[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel117_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel117 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111101010101100101011100110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel117[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel117_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel117 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111111001110110111111111111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel117[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel117_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel117 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b00111110101110101100010111101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel117[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel117_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel117 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111110010010101010011110010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel117[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel117_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel117 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111110000010111100100110011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel117[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel117_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel117 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111111011111000010110000100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel117[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel117_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel117 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111101110010000101010110110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel117[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel117_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel117 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b00111110100100000100001111100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel117[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel117_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel117 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b00111101010111110110100010111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel117[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel117_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel117 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111110111110000111000011011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel117[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel117_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel117 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111101110100111001010111001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel117[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel117_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel117 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111110001001100000010000100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel117[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel117_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel117 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b00111110010000110000111001001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel117[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel117_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel117 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111111000010100001100111110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel117[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel117_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel117 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111110111000010011000101001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel117[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel117_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel117 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111110000110111111101111110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel117[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel117_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel117 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111101011111101010100010010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel117[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel117_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel117 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111110110110010111101010101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel117[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel117_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel117 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b00111101100110010100011110011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel117[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel117_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel117 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111110001100111010001111000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel117[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel117_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel117 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111110100100101101101010110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel117[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel117_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel117 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111101001010101100111001001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel117[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel117_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel117 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111111000100101111010001010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel117[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel117_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel117 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b10111101010100001110011100110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel117[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel117_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel117 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111110101100011101001010111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel117[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel117_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel117 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111110100000111011100010100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel117[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel117_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel117 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111110011100111000101000101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel117[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel117_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel117 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111100100101110110001000001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel117[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel117_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel117 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111101100001101101111010010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel117[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel117_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel117 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111110100010010001110010110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel117[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel117_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel117 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b10111110110000011111011111010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel117[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel117_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel117 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b10111011000011010101001001001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel117[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel117_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel117 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111110100001010001100111001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel117[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel117_Valid_Out)
	);
	Adder_64input add_k117(
		.Data1(Data_Out_Kernel117[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel117[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel117[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel117[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel117[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel117[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel117[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel117[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel117[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel117[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel117[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel117[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel117[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel117[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel117[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel117[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel117[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel117[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel117[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel117[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel117[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel117[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel117[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel117[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel117[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel117[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel117[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel117[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel117[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel117[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel117[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel117[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel117[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel117[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel117[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel117[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel117[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel117[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel117[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel117[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel117[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel117[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel117[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel117[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel117[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel117[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel117[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel117[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel117[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel117[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel117[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel117[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel117[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel117[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel117[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel117[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel117[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel117[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel117[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel117[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel117[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel117[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel117[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel117[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel117),
		.Data_Out(add_k117_Data_Out),
		.Valid_Out(add_kernel117_Valid_Out)
	);
	Batch_Norm bn_kernel117(
		.Data_A(32'b00111101111111110010001100100101),
		.Data_B(32'b10111101000110111111100100110110),
		.Data_In(add_k117_Data_Out),
		.Valid_In(add_kernel117_Valid_Out),
		.Data_Out(bn117_Data_Out),
		.Valid_Out(bn117_Valid_Out)
	);
	Relu_Core rl_kernel117(
		.Data_In(bn117_Data_Out),
		.Valid_In(bn117_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*117-1:DATA_WIDHT*116]),
		.Valid_Out(rl117_Valid_Out)
	);
//////////KERNEL118//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel118 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110101111110101011011101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel118[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel118_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel118 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111101101100000101010101010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel118[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel118_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel118 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111100111011000111001100111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel118[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel118_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel118 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110100101100110001010011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel118[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel118_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel118 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111101010000010010001010101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel118[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel118_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel118 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110010000110010001000000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel118[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel118_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel118 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111110111001100100101011100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel118[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel118_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel118 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111111001110111010010101001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel118[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel118_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel118 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111110010011101011100101110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel118[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel118_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel118 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111111000000111111101100100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel118[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel118_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel118 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111111000101000011111010101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel118[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel118_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel118 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111110001011010110000001111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel118[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel118_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel118 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111111000100001011110111010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel118[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel118_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel118 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111110110000100111110001110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel118[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel118_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel118 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110100011111011001110110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel118[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel118_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel118 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111110100100110111010000111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel118[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel118_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel118 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111101000010111100001111011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel118[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel118_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel118 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111100111001010101100000001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel118[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel118_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel118 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111111000011111010001000101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel118[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel118_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel118 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111101111100000110101111001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel118[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel118_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel118 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111100110000110000001010010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel118[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel118_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel118 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111110100100011010001010011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel118[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel118_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel118 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110011001110111000001110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel118[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel118_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel118 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111110101001010100010001111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel118[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel118_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel118 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111101111101100010100011110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel118[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel118_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel118 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111101000011001010110110001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel118[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel118_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel118 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111111000000011110110001100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel118[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel118_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel118 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111111000101111111100101110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel118[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel118_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel118 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111110110010010101011011011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel118[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel118_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel118 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111111000000110110011010000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel118[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel118_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel118 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111110010110001111100000100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel118[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel118_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel118 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111111010111111010101110000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel118[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel118_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel118 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111110101111010010001110011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel118[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel118_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel118 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b00111110000000000111001010110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel118[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel118_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel118 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111110111010111000110111011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel118[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel118_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel118 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111101100111110011110001000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel118[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel118_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel118 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111110001101000001100100101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel118[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel118_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel118 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111111010001110101011010010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel118[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel118_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel118 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111111000110101001111001111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel118[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel118_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel118 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b00111110100011001001000011110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel118[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel118_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel118 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b10111110010110000101001001000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel118[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel118_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel118 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b10111110100110011001101110110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel118[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel118_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel118 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b00111101111001000011010010000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel118[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel118_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel118 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b00111101111001100001001110000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel118[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel118_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel118 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111110000010110001100001010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel118[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel118_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel118 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b10111110100101011100001110010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel118[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel118_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel118 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111110101010011010100101000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel118[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel118_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel118 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b00111110111011011111000010100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel118[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel118_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel118 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b00111110010001100000101000011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel118[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel118_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel118 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111110100100001001010011011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel118[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel118_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel118 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111110110000101100001011101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel118[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel118_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel118 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b10111110010001101001001011100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel118[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel118_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel118 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111110110000011100101100110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel118[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel118_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel118 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111101011011001100101100001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel118[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel118_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel118 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111110101010110111111011010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel118[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel118_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel118 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b00111111000101010100000010011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel118[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel118_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel118 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b10111101101010101101101101101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel118[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel118_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel118 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111110100110010011011010110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel118[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel118_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel118 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b10111110101100101101100100001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel118[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel118_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel118 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b00111111000010100100101110110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel118[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel118_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel118 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111110000011111111001101010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel118[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel118_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel118 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b10111110100111001101111100011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel118[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel118_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel118 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b10111101101101111000111000000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel118[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel118_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel118 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111101100011011101111011001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel118[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel118_Valid_Out)
	);
	Adder_64input add_k118(
		.Data1(Data_Out_Kernel118[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel118[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel118[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel118[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel118[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel118[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel118[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel118[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel118[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel118[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel118[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel118[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel118[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel118[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel118[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel118[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel118[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel118[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel118[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel118[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel118[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel118[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel118[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel118[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel118[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel118[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel118[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel118[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel118[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel118[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel118[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel118[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel118[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel118[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel118[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel118[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel118[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel118[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel118[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel118[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel118[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel118[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel118[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel118[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel118[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel118[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel118[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel118[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel118[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel118[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel118[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel118[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel118[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel118[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel118[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel118[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel118[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel118[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel118[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel118[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel118[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel118[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel118[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel118[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel118),
		.Data_Out(add_k118_Data_Out),
		.Valid_Out(add_kernel118_Valid_Out)
	);
	Batch_Norm bn_kernel118(
		.Data_A(32'b00111110001111011010111110001110),
		.Data_B(32'b00111111100010110100100001111100),
		.Data_In(add_k118_Data_Out),
		.Valid_In(add_kernel118_Valid_Out),
		.Data_Out(bn118_Data_Out),
		.Valid_Out(bn118_Valid_Out)
	);
	Relu_Core rl_kernel118(
		.Data_In(bn118_Data_Out),
		.Valid_In(bn118_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*118-1:DATA_WIDHT*117]),
		.Valid_Out(rl118_Valid_Out)
	);
//////////KERNEL119//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel119 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111111000100101100110101100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel119[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel119_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel119 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110000100001101101011100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel119[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel119_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel119 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110000010100000001100001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel119[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel119_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel119 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110100100111000111010001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel119[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel119_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel119 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111101111001110000111111001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel119[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel119_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel119 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111101100100110101000011110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel119[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel119_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel119 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111110001010000001001011010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel119[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel119_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel119 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111110001011110000010100101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel119[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel119_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel119 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110100100101011111100011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel119[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel119_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel119 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111100100100100111111101011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel119[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel119_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel119 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111110011000001000010010011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel119[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel119_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel119 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111110101001011101010101111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel119[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel119_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel119 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110001011111111010001111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel119[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel119_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel119 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111101100101010110100110111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel119[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel119_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel119 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110100111111010100001011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel119[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel119_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel119 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111101001010110111110010111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel119[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel119_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel119 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110101111110110010010110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel119[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel119_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel119 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111101100010001000001000100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel119[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel119_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel119 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110110011001110101101110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel119[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel119_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel119 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110011111010000100011011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel119[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel119_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel119 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110001001100000101001101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel119[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel119_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel119 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111101001010011111011111110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel119[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel119_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel119 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110111001011101010110100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel119[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel119_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel119 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111110000111100011101011100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel119[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel119_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel119 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111101100001110001001110111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel119[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel119_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel119 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110010011100101101100111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel119[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel119_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel119 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110001100001111100000100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel119[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel119_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel119 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111101101101101010000000011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel119[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel119_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel119 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111101100100000110010011001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel119[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel119_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel119 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111110101111101101111000101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel119[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel119_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel119 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111101000101011100110110100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel119[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel119_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel119 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111100110001010110111100000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel119[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel119_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel119 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b00111110010100110010001100001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel119[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel119_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel119 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b00111101100000000111010111010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel119[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel119_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel119 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111110110101001110010010010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel119[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel119_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel119 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b10111100100001110101111011100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel119[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel119_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel119 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111110110000010100110011100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel119[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel119_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel119 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111011101010101110101100100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel119[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel119_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel119 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b00111101110101111100101101011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel119[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel119_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel119 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111101011010010000011001101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel119[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel119_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel119 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111111000110000000100110100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel119[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel119_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel119 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111101011010110011010100011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel119[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel119_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel119 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111110001101101111011011100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel119[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel119_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel119 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111110101010001111000011001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel119[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel119_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel119 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111101001010000010110101111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel119[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel119_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel119 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111110010101110001001010110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel119[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel119_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel119 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111110101101001111111011001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel119[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel119_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel119 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111110100011000000010000001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel119[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel119_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel119 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111110000111001010111000010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel119[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel119_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel119 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111110000110111010011001000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel119[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel119_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel119 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111110001101011001000111100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel119[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel119_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel119 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111100001100001000111100111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel119[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel119_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel119 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111110010000001100111100111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel119[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel119_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel119 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111110100001001000010011010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel119[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel119_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel119 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111101010111011010000011111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel119[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel119_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel119 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b00111110001010110010101111001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel119[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel119_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel119 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111110011101111010101000111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel119[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel119_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel119 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111110000010010001001111010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel119[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel119_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel119 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b10111100100011100010001000000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel119[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel119_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel119 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b00111101001110100010111101010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel119[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel119_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel119 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111110001101000100000101001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel119[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel119_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel119 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b10111100111001111001111000111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel119[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel119_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel119 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111110001010011100000001110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel119[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel119_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel119 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b10111101010010110011011101100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel119[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel119_Valid_Out)
	);
	Adder_64input add_k119(
		.Data1(Data_Out_Kernel119[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel119[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel119[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel119[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel119[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel119[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel119[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel119[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel119[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel119[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel119[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel119[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel119[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel119[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel119[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel119[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel119[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel119[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel119[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel119[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel119[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel119[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel119[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel119[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel119[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel119[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel119[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel119[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel119[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel119[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel119[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel119[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel119[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel119[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel119[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel119[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel119[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel119[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel119[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel119[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel119[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel119[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel119[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel119[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel119[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel119[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel119[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel119[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel119[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel119[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel119[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel119[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel119[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel119[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel119[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel119[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel119[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel119[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel119[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel119[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel119[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel119[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel119[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel119[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel119),
		.Data_Out(add_k119_Data_Out),
		.Valid_Out(add_kernel119_Valid_Out)
	);
	Batch_Norm bn_kernel119(
		.Data_A(32'b00111110011101001111010111111011),
		.Data_B(32'b10111110101101111001010000000100),
		.Data_In(add_k119_Data_Out),
		.Valid_In(add_kernel119_Valid_Out),
		.Data_Out(bn119_Data_Out),
		.Valid_Out(bn119_Valid_Out)
	);
	Relu_Core rl_kernel119(
		.Data_In(bn119_Data_Out),
		.Valid_In(bn119_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*119-1:DATA_WIDHT*118]),
		.Valid_Out(rl119_Valid_Out)
	);
//////////KERNEL120//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel120 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110100011010000010101000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel120[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel120_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel120 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111101111011001101001010000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel120[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel120_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel120 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111111001111110000001001101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel120[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel120_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel120 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110111011101110110001010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel120[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel120_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel120 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111110011110110110100000010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel120[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel120_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel120 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111100110100010101110010001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel120[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel120_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel120 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111111001001101011101101111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel120[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel120_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel120 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111111001001101110111000010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel120[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel120_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel120 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111111001011100100011010000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel120[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel120_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel120 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110010000111110101100111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel120[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel120_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel120 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111101010111001001110010100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel120[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel120_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel120 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111101100111001111010001101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel120[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel120_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel120 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110110111110101110101010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel120[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel120_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel120 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111110011100100110011001100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel120[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel120_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel120 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110010010011010111001110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel120[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel120_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel120 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111111001001110011100111001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel120[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel120_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel120 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111110100100010110010101100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel120[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel120_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel120 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110001011010101111000000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel120[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel120_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel120 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111101001111110111110111000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel120[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel120_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel120 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110100111100010101010101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel120[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel120_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel120 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111101100111000101010110000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel120[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel120_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel120 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111110001100000100101110100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel120[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel120_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel120 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110000111100110110101001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel120[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel120_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel120 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111111010011011000011101001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel120[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel120_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel120 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111110110111001010110101100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel120[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel120_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel120 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111111000010000010110100011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel120[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel120_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel120 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111101100001011100011000001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel120[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel120_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel120 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111111000011110000100010101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel120[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel120_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel120 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111110111100100110010010111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel120[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel120_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel120 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110010001110101001110011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel120[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel120_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel120 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111100001101001011000010110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel120[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel120_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel120 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111101001100110110000101100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel120[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel120_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel120 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111101010101100010011000000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel120[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel120_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel120 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b00111101110000111000110011101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel120[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel120_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel120 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111110100010001111101011010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel120[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel120_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel120 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b10111100101110010110111101101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel120[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel120_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel120 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b10111110000110110000010010100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel120[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel120_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel120 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111110011000010000110110011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel120[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel120_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel120 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111111001000001001000100111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel120[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel120_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel120 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111110000110111110000110001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel120[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel120_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel120 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b10111110101000111010001011011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel120[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel120_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel120 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111110000110100011001110000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel120[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel120_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel120 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b00111101110101000011011100000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel120[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel120_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel120 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b00111110000001001110000001011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel120[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel120_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel120 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111110011010101111011101111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel120[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel120_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel120 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b10111111010000110001100110101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel120[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel120_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel120 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b10111101100011100101110011110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel120[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel120_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel120 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b00111110001111001110110111111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel120[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel120_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel120 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111101010010111101001111111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel120[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel120_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel120 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b00111110001100000110110101110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel120[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel120_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel120 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111110010001001001101001110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel120[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel120_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel120 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b10111110010011011110100001011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel120[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel120_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel120 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111110100001101010001010100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel120[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel120_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel120 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b00111110101010000100011000110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel120[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel120_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel120 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111110001010011011001100111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel120[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel120_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel120 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b00111111001101110100110101001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel120[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel120_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel120 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b10111111001000101000111010101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel120[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel120_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel120 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b10111100010000100111110111100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel120[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel120_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel120 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b10111110011100001000111100100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel120[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel120_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel120 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111111000001000011101100010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel120[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel120_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel120 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111110001100010000101110111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel120[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel120_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel120 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b10111101001011000110111001100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel120[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel120_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel120 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111101010001101100010001100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel120[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel120_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel120 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b10111101111000000101000010011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel120[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel120_Valid_Out)
	);
	Adder_64input add_k120(
		.Data1(Data_Out_Kernel120[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel120[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel120[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel120[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel120[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel120[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel120[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel120[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel120[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel120[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel120[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel120[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel120[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel120[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel120[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel120[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel120[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel120[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel120[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel120[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel120[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel120[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel120[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel120[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel120[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel120[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel120[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel120[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel120[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel120[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel120[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel120[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel120[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel120[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel120[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel120[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel120[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel120[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel120[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel120[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel120[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel120[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel120[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel120[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel120[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel120[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel120[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel120[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel120[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel120[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel120[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel120[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel120[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel120[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel120[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel120[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel120[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel120[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel120[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel120[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel120[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel120[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel120[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel120[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel120),
		.Data_Out(add_k120_Data_Out),
		.Valid_Out(add_kernel120_Valid_Out)
	);
	Batch_Norm bn_kernel120(
		.Data_A(32'b00111110000101101111011011100111),
		.Data_B(32'b00111111001110110111000010111010),
		.Data_In(add_k120_Data_Out),
		.Valid_In(add_kernel120_Valid_Out),
		.Data_Out(bn120_Data_Out),
		.Valid_Out(bn120_Valid_Out)
	);
	Relu_Core rl_kernel120(
		.Data_In(bn120_Data_Out),
		.Valid_In(bn120_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*120-1:DATA_WIDHT*119]),
		.Valid_Out(rl120_Valid_Out)
	);
//////////KERNEL121//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel121 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111101111011111001111101111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel121[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel121_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel121 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110100000111110111011010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel121[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel121_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel121 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110110011000100110101110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel121[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel121_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel121 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110101110000100111111101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel121[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel121_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel121 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111110001101011110110101010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel121[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel121_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel121 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110010001001000011000000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel121[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel121_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel121 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111111001011001010011001101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel121[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel121_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel121 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111110001001011001100010101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel121[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel121_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel121 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111111001011011000111000100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel121[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel121_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel121 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111101100001000011101100010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel121[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel121_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel121 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110001010001001101110110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel121[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel121_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel121 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111110010111100100011100000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel121[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel121_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel121 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111101101101101100101011010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel121[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel121_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel121 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111110001011100110001100001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel121[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel121_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel121 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111101100110111000100001001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel121[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel121_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel121 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111110100000100110010000110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel121[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel121_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel121 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110110000001110000000111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel121[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel121_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel121 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111110100101011100101100000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel121[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel121_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel121 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111111000100010010001110110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel121[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel121_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel121 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111100110101110100010100010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel121[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel121_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel121 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111111000011111000110111011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel121[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel121_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel121 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111110100111001010110010000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel121[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel121_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel121 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110111100011110000110110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel121[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel121_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel121 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111111010111100110100011011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel121[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel121_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel121 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111101110001100000110010011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel121[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel121_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel121 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111101000101111011111110101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel121[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel121_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel121 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111111000000010100010011100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel121[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel121_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel121 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110011001110110001010000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel121[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel121_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel121 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111110111100000111101100000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel121[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel121_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel121 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110011111100101001010011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel121[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel121_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel121 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111111000001110110111001000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel121[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel121_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel121 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110111001110100000100011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel121[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel121_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel121 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111110101101000011001101100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel121[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel121_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel121 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b00111111000101010001010000001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel121[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel121_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel121 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111110110110111101110101000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel121[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel121_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel121 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b10111101000000011001011010111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel121[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel121_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel121 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111111001100001011001100101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel121[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel121_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel121 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111110010001100000010000110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel121[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel121_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel121 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b00111101110100110000100001111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel121[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel121_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel121 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111100011110011001110011010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel121[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel121_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel121 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111111000101001111000101001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel121[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel121_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel121 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b10111110000101111000110101001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel121[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel121_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel121 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111101101100110011101100111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel121[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel121_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel121 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111101101010101001111000101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel121[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel121_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel121 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111110100010001001000110101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel121[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel121_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel121 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111110110001111000000001001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel121[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel121_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel121 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111110000010110100000110101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel121[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel121_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel121 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111110010110000101001101100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel121[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel121_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel121 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111110101011001011110101110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel121[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel121_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel121 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b00111110000010000101101010001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel121[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel121_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel121 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111100000100000001001110100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel121[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel121_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel121 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111110011000010100111100011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel121[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel121_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel121 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b00111110101010000000101011001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel121[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel121_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel121 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111110101001110110001101001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel121[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel121_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel121 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b10111101110101010100101010111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel121[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel121_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel121 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111111001010000011101001010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel121[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel121_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel121 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111110000010101101110111110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel121[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel121_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel121 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b10111101111011110000110100001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel121[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel121_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel121 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b10111110010110011110011111000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel121[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel121_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel121 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b00111110001100100010100111010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel121[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel121_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel121 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b10111110011001100011010001011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel121[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel121_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel121 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b10111011111110010011111011111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel121[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel121_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel121 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b10111101101010010011010000101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel121[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel121_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel121 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111110000110000101101001110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel121[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel121_Valid_Out)
	);
	Adder_64input add_k121(
		.Data1(Data_Out_Kernel121[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel121[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel121[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel121[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel121[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel121[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel121[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel121[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel121[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel121[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel121[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel121[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel121[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel121[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel121[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel121[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel121[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel121[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel121[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel121[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel121[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel121[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel121[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel121[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel121[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel121[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel121[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel121[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel121[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel121[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel121[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel121[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel121[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel121[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel121[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel121[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel121[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel121[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel121[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel121[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel121[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel121[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel121[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel121[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel121[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel121[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel121[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel121[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel121[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel121[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel121[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel121[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel121[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel121[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel121[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel121[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel121[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel121[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel121[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel121[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel121[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel121[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel121[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel121[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel121),
		.Data_Out(add_k121_Data_Out),
		.Valid_Out(add_kernel121_Valid_Out)
	);
	Batch_Norm bn_kernel121(
		.Data_A(32'b00111110000000100110111110010000),
		.Data_B(32'b10111110000001011101100010000001),
		.Data_In(add_k121_Data_Out),
		.Valid_In(add_kernel121_Valid_Out),
		.Data_Out(bn121_Data_Out),
		.Valid_Out(bn121_Valid_Out)
	);
	Relu_Core rl_kernel121(
		.Data_In(bn121_Data_Out),
		.Valid_In(bn121_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*121-1:DATA_WIDHT*120]),
		.Valid_Out(rl121_Valid_Out)
	);
//////////KERNEL122//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel122 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111110100011011000110100100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel122[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel122_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel122 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110001001001111000100011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel122[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel122_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel122 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110100100001010111111011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel122[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel122_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel122 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110100100100101110000010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel122[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel122_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel122 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111100101101111110011001101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel122[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel122_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel122 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111101101110010110101011101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel122[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel122_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel122 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111110001111010010010000000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel122[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel122_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel122 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111101100100111111000111111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel122[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel122_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel122 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111101001010000000100111011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel122[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel122_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel122 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111110100000001010100000101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel122[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel122_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel122 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111100111111001111110110000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel122[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel122_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel122 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111100101011100100110111010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel122[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel122_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel122 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110000011000110010001110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel122[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel122_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel122 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111101111010110001000100111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel122[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel122_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel122 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111101111011100000001000000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel122[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel122_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel122 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111101100001110100111111000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel122[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel122_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel122 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110011010111000101001111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel122[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel122_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel122 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111101101111010010101111110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel122[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel122_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel122 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111101100101100101010110001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel122[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel122_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel122 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110110011010010101100001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel122[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel122_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel122 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110110011000110110101100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel122[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel122_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel122 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111110100011111001110101011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel122[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel122_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel122 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111101100001001000110100001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel122[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel122_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel122 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111110100101001001101111001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel122[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel122_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel122 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111100110101001010000001110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel122[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel122_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel122 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110100110011011001100100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel122[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel122_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel122 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110101100111001110101101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel122[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel122_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel122 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110111000110010001000000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel122[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel122_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel122 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111110001100110010001000100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel122[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel122_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel122 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111101101100010011111110111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel122[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel122_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel122 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111110011110101000011011110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel122[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel122_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel122 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110010001001100100011101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel122[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel122_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel122 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111110111000111100110100101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel122[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel122_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel122 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b00111110111001010110111100011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel122[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel122_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel122 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111111001001110110101010100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel122[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel122_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel122 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b10111110000000010100111001000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel122[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel122_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel122 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111110001100001011100100011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel122[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel122_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel122 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111101111010011100010101110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel122[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel122_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel122 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b00111101101111101110101000010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel122[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel122_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel122 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b00111100011011110000010000000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel122[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel122_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel122 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111111000000011001110101110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel122[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel122_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel122 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111110010001100001100111100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel122[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel122_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel122 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b00111110000100011101110000101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel122[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel122_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel122 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b00111100101110100010010000110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel122[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel122_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel122 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111110110111011001100110011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel122[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel122_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel122 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111110101100111100111010100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel122[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel122_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel122 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111101011101011101001000000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel122[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel122_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel122 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111111000111101000111001011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel122[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel122_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel122 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111101101110001101000100010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel122[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel122_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel122 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b00111101010101101100110111000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel122[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel122_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel122 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111101000111110010001010011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel122[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel122_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel122 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111110111101111001000110000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel122[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel122_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel122 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b00111110101001110111100111001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel122[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel122_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel122 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111111000111100101110001011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel122[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel122_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel122 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111011000100111011101110100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel122[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel122_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel122 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111110100110011000110101100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel122[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel122_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel122 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111110110101100100111101001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel122[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel122_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel122 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111101000011111100000010000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel122[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel122_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel122 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b10111110100100110110101000001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel122[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel122_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel122 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b00111110100111011000011111011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel122[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel122_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel122 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111101011111100010100000111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel122[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel122_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel122 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b10111110011000110001001111100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel122[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel122_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel122 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b10111100111111100101000100001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel122[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel122_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel122 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b10111101100001000110010001100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel122[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel122_Valid_Out)
	);
	Adder_64input add_k122(
		.Data1(Data_Out_Kernel122[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel122[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel122[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel122[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel122[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel122[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel122[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel122[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel122[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel122[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel122[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel122[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel122[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel122[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel122[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel122[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel122[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel122[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel122[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel122[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel122[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel122[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel122[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel122[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel122[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel122[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel122[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel122[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel122[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel122[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel122[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel122[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel122[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel122[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel122[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel122[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel122[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel122[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel122[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel122[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel122[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel122[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel122[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel122[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel122[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel122[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel122[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel122[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel122[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel122[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel122[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel122[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel122[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel122[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel122[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel122[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel122[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel122[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel122[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel122[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel122[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel122[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel122[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel122[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel122),
		.Data_Out(add_k122_Data_Out),
		.Valid_Out(add_kernel122_Valid_Out)
	);
	Batch_Norm bn_kernel122(
		.Data_A(32'b00111110001111100110101000110100),
		.Data_B(32'b10111110111101100100110101101100),
		.Data_In(add_k122_Data_Out),
		.Valid_In(add_kernel122_Valid_Out),
		.Data_Out(bn122_Data_Out),
		.Valid_Out(bn122_Valid_Out)
	);
	Relu_Core rl_kernel122(
		.Data_In(bn122_Data_Out),
		.Valid_In(bn122_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*122-1:DATA_WIDHT*121]),
		.Valid_Out(rl122_Valid_Out)
	);
//////////KERNEL123//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel123 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110010001100001101101001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel123[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel123_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel123 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111110001100100111011001000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel123[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel123_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel123 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110010101100110111000100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel123[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel123_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel123 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110101110110100011111111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel123[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel123_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel123 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111101000101101010001100001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel123[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel123_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel123 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111101010010111101011100101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel123[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel123_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel123 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111110100010010010010001010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel123[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel123_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel123 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111100101111010101000010100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel123[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel123_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel123 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111110100010000111001111011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel123[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel123_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel123 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110000101110011010000010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel123[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel123_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel123 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111101101010011000100001011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel123[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel123_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel123 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111010110110000010011110001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel123[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel123_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel123 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110000100110101010011100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel123[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel123_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel123 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111110101101000110011100100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel123[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel123_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel123 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110100111000001000001111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel123[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel123_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel123 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111110100101100111101011001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel123[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel123_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel123 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111101001000111000010110011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel123[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel123_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel123 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111101111111011110000001100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel123[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel123_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel123 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111101100010011010010011010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel123[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel123_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel123 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111101010101000110111010011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel123[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel123_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel123 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110101111011001100100100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel123[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel123_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel123 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111101111001110010110110100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel123[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel123_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel123 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111110100011011010001111001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel123[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel123_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel123 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111110100111101011011101100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel123[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel123_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel123 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111101000000101100001101011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel123[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel123_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel123 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111110011000011000101001010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel123[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel123_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel123 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111110111000000110001100001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel123[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel123_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel123 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111110111111011111010101111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel123[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel123_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel123 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111110000100001100111100111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel123[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel123_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel123 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111111000100100110100111101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel123[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel123_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel123 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111110001101000010100110110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel123[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel123_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel123 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111100000100011100100010110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel123[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel123_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel123 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b00111110001101101010111111010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel123[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel123_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel123 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111110111011110000001110000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel123[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel123_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel123 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111111010101100110010101110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel123[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel123_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel123 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111110010100000100110010110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel123[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel123_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel123 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111011100111111111111000100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel123[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel123_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel123 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b00111101101011000110011010001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel123[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel123_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel123 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111110101011100100000111110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel123[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel123_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel123 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111100100110100000000101111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel123[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel123_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel123 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b10111110101101110100111111110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel123[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel123_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel123 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111110001011111101100110111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel123[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel123_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel123 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b00111101000011100011000000001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel123[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel123_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel123 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b10111100100001110111111111010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel123[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel123_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel123 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b00111110101001010001111001000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel123[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel123_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel123 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b10111110100001111100110011011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel123[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel123_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel123 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111101011010111110100101010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel123[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel123_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel123 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b00111110111000100010010011011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel123[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel123_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel123 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b00111101111101001010111010110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel123[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel123_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel123 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b00111110011001011110001011001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel123[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel123_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel123 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111101010101010101000111101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel123[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel123_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel123 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b10111110111000111010100101001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel123[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel123_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel123 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111110011110100110110001100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel123[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel123_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel123 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b00111110100011010011011000001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel123[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel123_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel123 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b10111101100000000000011011001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel123[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel123_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel123 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b00111110011001001101001001100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel123[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel123_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel123 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b10111110110111101010110110101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel123[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel123_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel123 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b10111110100100111111110111111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel123[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel123_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel123 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111110011111100110001001100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel123[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel123_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel123 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b00111101000101011001110100001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel123[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel123_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel123 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111110001100010000011110101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel123[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel123_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel123 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111110000101001101111110010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel123[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel123_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel123 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b10111101101001010101111111010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel123[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel123_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel123 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111110000010011001000101101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel123[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel123_Valid_Out)
	);
	Adder_64input add_k123(
		.Data1(Data_Out_Kernel123[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel123[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel123[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel123[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel123[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel123[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel123[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel123[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel123[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel123[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel123[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel123[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel123[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel123[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel123[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel123[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel123[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel123[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel123[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel123[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel123[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel123[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel123[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel123[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel123[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel123[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel123[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel123[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel123[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel123[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel123[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel123[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel123[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel123[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel123[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel123[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel123[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel123[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel123[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel123[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel123[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel123[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel123[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel123[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel123[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel123[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel123[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel123[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel123[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel123[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel123[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel123[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel123[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel123[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel123[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel123[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel123[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel123[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel123[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel123[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel123[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel123[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel123[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel123[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel123),
		.Data_Out(add_k123_Data_Out),
		.Valid_Out(add_kernel123_Valid_Out)
	);
	Batch_Norm bn_kernel123(
		.Data_A(32'b00111110010001011011100100000010),
		.Data_B(32'b10111101101101110011000100100101),
		.Data_In(add_k123_Data_Out),
		.Valid_In(add_kernel123_Valid_Out),
		.Data_Out(bn123_Data_Out),
		.Valid_Out(bn123_Valid_Out)
	);
	Relu_Core rl_kernel123(
		.Data_In(bn123_Data_Out),
		.Valid_In(bn123_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*123-1:DATA_WIDHT*122]),
		.Valid_Out(rl123_Valid_Out)
	);
//////////KERNEL124//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel124 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111110101101110101010011010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel124[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel124_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel124 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111101110011010100111011101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel124[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel124_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel124 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110101011110100110101111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel124[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel124_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel124 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110101111111001001111001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel124[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel124_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel124 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111101011101111110001010010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel124[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel124_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel124 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110100101101100010111010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel124[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel124_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel124 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111110001111100000100000101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel124[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel124_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel124 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111101110000110101101101110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel124[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel124_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel124 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111101010101000101101101101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel124[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel124_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel124 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111100111001001101011101001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel124[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel124_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel124 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111100111001000000010100101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel124[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel124_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel124 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111101100100111011110101111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel124[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel124_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel124 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111101111000110110111010100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel124[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel124_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel124 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111110001000111101111100101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel124[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel124_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel124 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110001110100111111010001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel124[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel124_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel124 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111110001010101100001111111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel124[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel124_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel124 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110001100101111101111011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel124[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel124_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel124 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110001000100011111101010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel124[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel124_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel124 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111101011011000101010001011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel124[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel124_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel124 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111101010001100011000000100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel124[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel124_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel124 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110100110011011000000100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel124[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel124_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel124 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111101101010111001101111100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel124[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel124_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel124 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111111001110101001100110100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel124[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel124_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel124 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111110010011010010011100110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel124[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel124_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel124 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111110011101010011001010100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel124[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel124_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel124 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110010001111100101010111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel124[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel124_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel124 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110011111010101001101110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel124[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel124_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel124 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110100001011001000110100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel124[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel124_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel124 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111110100000000101011011010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel124[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel124_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel124 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111110101000101111010111010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel124[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel124_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel124 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111110100111010010111010110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel124[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel124_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel124 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110011011101010001010000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel124[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel124_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel124 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111111001001111101001101001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel124[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel124_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel124 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b00111110001001000011011000000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel124[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel124_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel124 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111111001001111011100011000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel124[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel124_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel124 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b10111110100010110110100001001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel124[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel124_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel124 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111110110100110101011101001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel124[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel124_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel124 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111110000000111110100000100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel124[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel124_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel124 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b00111110010011101011100011110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel124[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel124_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel124 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111110011110001010111011011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel124[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel124_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel124 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111111000110100001010111100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel124[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel124_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel124 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111110011100000001010110111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel124[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel124_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel124 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111110000111000101011001101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel124[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel124_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel124 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b00111101110100001101110010110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel124[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel124_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel124 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111111000100001110000110101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel124[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel124_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel124 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111110100101010010000100011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel124[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel124_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel124 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111110001110001100101110000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel124[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel124_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel124 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111101100111111010010100110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel124[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel124_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel124 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111110011111100101100110101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel124[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel124_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel124 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b00111100111010101010011010111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel124[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel124_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel124 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111110111001111000000010110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel124[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel124_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel124 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111110100100011110110000010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel124[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel124_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel124 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b00111101101111011111000010010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel124[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel124_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel124 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111111001010111000110100011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel124[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel124_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel124 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111110101110111110011110100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel124[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel124_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel124 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111110010000001111000101101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel124[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel124_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel124 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111110011011010111000111000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel124[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel124_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel124 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111110010000011110100111111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel124[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel124_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel124 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111101110001110101000001011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel124[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel124_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel124 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111101110010100110010101110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel124[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel124_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel124 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111110111100000101011101111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel124[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel124_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel124 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111100101010011100010101001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel124[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel124_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel124 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111110011111110111100000101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel124[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel124_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel124 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111101110000010100001010010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel124[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel124_Valid_Out)
	);
	Adder_64input add_k124(
		.Data1(Data_Out_Kernel124[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel124[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel124[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel124[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel124[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel124[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel124[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel124[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel124[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel124[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel124[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel124[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel124[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel124[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel124[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel124[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel124[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel124[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel124[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel124[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel124[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel124[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel124[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel124[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel124[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel124[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel124[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel124[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel124[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel124[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel124[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel124[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel124[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel124[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel124[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel124[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel124[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel124[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel124[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel124[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel124[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel124[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel124[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel124[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel124[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel124[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel124[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel124[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel124[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel124[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel124[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel124[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel124[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel124[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel124[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel124[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel124[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel124[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel124[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel124[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel124[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel124[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel124[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel124[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel124),
		.Data_Out(add_k124_Data_Out),
		.Valid_Out(add_kernel124_Valid_Out)
	);
	Batch_Norm bn_kernel124(
		.Data_A(32'b00111110001010011001010100000110),
		.Data_B(32'b10111110110101110011000010011101),
		.Data_In(add_k124_Data_Out),
		.Valid_In(add_kernel124_Valid_Out),
		.Data_Out(bn124_Data_Out),
		.Valid_Out(bn124_Valid_Out)
	);
	Relu_Core rl_kernel124(
		.Data_In(bn124_Data_Out),
		.Valid_In(bn124_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*124-1:DATA_WIDHT*123]),
		.Valid_Out(rl124_Valid_Out)
	);
//////////KERNEL125//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel125 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110110011010000010000111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel125[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel125_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel125 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111110101110010110100010100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel125[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel125_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel125 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111101101011001000111111010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel125[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel125_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel125 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110100000010100001110100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel125[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel125_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel125 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111110001101001100110100001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel125[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel125_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel125 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111101000111010010101110011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel125[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel125_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel125 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111110001111010001000100000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel125[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel125_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel125 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111110001010111110101100110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel125[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel125_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel125 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111110110010011111110001001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel125[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel125_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel125 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110011001100001110000000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel125[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel125_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel125 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111101111100010010111010101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel125[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel125_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel125 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110001101111000100111011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel125[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel125_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel125 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111101100100100001011001110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel125[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel125_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel125 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111110100000001100001111100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel125[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel125_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel125 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110110001111000100011011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel125[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel125_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel125 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111100110101000110000000101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel125[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel125_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel125 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111101110011111111010011111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel125[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel125_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel125 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111101111011001110010110111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel125[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel125_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel125 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111100101001001011011110010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel125[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel125_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel125 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111100110100111100100100001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel125[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel125_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel125 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110110000011000011011000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel125[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel125_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel125 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111100011101010110101110011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel125[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel125_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel125 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111111000011100011100111011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel125[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel125_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel125 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111101111110110110000010001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel125[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel125_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel125 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111101101000100011001100100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel125[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel125_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel125 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111101110010011100010111110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel125[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel125_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel125 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111110110101100010110010100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel125[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel125_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel125 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111111000100110000000000000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel125[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel125_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel125 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111101010110001101111011100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel125[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel125_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel125 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110111110001000100010010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel125[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel125_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel125 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111110001011001101101110011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel125[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel125_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel125 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111110001000101101001001000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel125[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel125_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel125 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b00111110000010111110001111011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel125[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel125_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel125 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111110110111110000111000111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel125[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel125_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel125 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111111000101100000001010101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel125[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel125_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel125 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111110000010001001101010001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel125[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel125_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel125 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b10111110010111100110101001100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel125[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel125_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel125 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b10111100101001101111111011111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel125[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel125_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel125 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111110100000011101110111111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel125[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel125_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel125 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111101101111101101111110101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel125[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel125_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel125 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b10111111000001110001100011001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel125[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel125_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel125 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111011100111110001100101110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel125[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel125_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel125 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b00111110011011010101000000001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel125[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel125_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel125 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b00111101101001110101011100011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel125[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel125_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel125 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b00111110100101011011000010001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel125[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel125_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel125 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b10111110000111000100110000110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel125[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel125_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel125 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b10111110010001100000010111111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel125[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel125_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel125 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b00111110101110011110100011011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel125[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel125_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel125 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b00111100111011100000111111000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel125[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel125_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel125 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b00111110000010111000011010110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel125[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel125_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel125 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111101101111010011101111110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel125[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel125_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel125 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b10111110000110010111110001101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel125[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel125_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel125 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111101100110000100010101001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel125[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel125_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel125 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b00111101101000001010111101011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel125[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel125_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel125 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b10111101101101111110001000000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel125[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel125_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel125 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b00111100100110110001101111111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel125[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel125_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel125 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b10111110011001011100011011001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel125[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel125_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel125 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b10111110111011101110100100001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel125[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel125_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel125 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111110111010100001101101011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel125[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel125_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel125 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111100010011111010110101010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel125[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel125_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel125 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b10111101110101001111001100100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel125[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel125_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel125 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111101011110001011111111101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel125[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel125_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel125 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b10111101110111111010100001101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel125[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel125_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel125 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111110011001110010001101001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel125[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel125_Valid_Out)
	);
	Adder_64input add_k125(
		.Data1(Data_Out_Kernel125[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel125[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel125[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel125[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel125[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel125[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel125[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel125[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel125[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel125[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel125[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel125[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel125[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel125[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel125[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel125[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel125[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel125[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel125[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel125[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel125[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel125[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel125[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel125[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel125[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel125[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel125[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel125[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel125[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel125[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel125[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel125[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel125[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel125[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel125[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel125[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel125[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel125[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel125[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel125[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel125[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel125[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel125[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel125[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel125[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel125[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel125[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel125[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel125[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel125[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel125[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel125[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel125[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel125[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel125[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel125[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel125[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel125[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel125[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel125[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel125[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel125[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel125[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel125[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel125),
		.Data_Out(add_k125_Data_Out),
		.Valid_Out(add_kernel125_Valid_Out)
	);
	Batch_Norm bn_kernel125(
		.Data_A(32'b00111110010100101110010001000001),
		.Data_B(32'b10111101011011011010001000011111),
		.Data_In(add_k125_Data_Out),
		.Valid_In(add_kernel125_Valid_Out),
		.Data_Out(bn125_Data_Out),
		.Valid_Out(bn125_Valid_Out)
	);
	Relu_Core rl_kernel125(
		.Data_In(bn125_Data_Out),
		.Valid_In(bn125_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*125-1:DATA_WIDHT*124]),
		.Valid_Out(rl125_Valid_Out)
	);
//////////KERNEL126//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel126 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110101001000010010111000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel126[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel126_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel126 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111110110100111110110001100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel126[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel126_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel126 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110101100101001100111101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel126[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel126_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel126 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110110010111000000001000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel126[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel126_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel126 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111101110111110000001111101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel126[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel126_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel126 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111100110100100011110000001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel126[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel126_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel126 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111110101101110000110101100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel126[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel126_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel126 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111101011101110001100111011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel126[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel126_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel126 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111101110100010100011101011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel126[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel126_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel126 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111101100000101101010011110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel126[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel126_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel126 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111011011011000111010100100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel126[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel126_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel126 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110001010010101100010011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel126[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel126_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel126 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110000010110101100100100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel126[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel126_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel126 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111110000000011001000111000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel126[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel126_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel126 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110111000111001101111010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel126[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel126_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel126 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111110010110010010111001000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel126[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel126_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel126 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111110101111110000001000101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel126[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel126_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel126 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111110100100000101001100010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel126[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel126_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel126 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111101101000110111101100010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel126[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel126_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel126 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111101100011010001001100100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel126[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel126_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel126 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110000010100011101011111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel126[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel126_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel126 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111101101011110100100010000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel126[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel126_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel126 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111101110100110111100110001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel126[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel126_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel126 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111110011011001001110100000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel126[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel126_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel126 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111101010100000000001110101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel126[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel126_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel126 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111101111110010100010110000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel126[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel126_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel126 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111110111100111001011100101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel126[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel126_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel126 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111110100100111000100011100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel126[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel126_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel126 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111110001011000101010011010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel126[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel126_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel126 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110111100010100101110101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel126[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel126_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel126 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111110011100010100101010101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel126[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel126_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel126 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111110110000001111111100110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel126[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel126_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel126 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111110001001000100100011011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel126[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel126_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel126 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111110010000011010101101000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel126[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel126_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel126 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b10111110101101110010111101111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel126[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel126_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel126 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111101101001010011110111001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel126[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel126_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel126 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b10111101001110110010100111010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel126[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel126_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel126 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b00111101110100010110111010001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel126[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel126_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel126 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b10111110011100001000010001100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel126[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel126_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel126 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b00111101110001001101110001000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel126[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel126_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel126 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b10111111010001010100011110100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel126[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel126_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel126 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111100111010001110010011001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel126[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel126_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel126 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b00111101110011100101111001110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel126[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel126_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel126 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b00111110100000100001001001100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel126[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel126_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel126 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b00111110011011111100100111011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel126[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel126_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel126 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b10111110010011000011100010011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel126[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel126_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel126 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b10111110000111101111001010000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel126[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel126_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel126 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b00111110101000100011010010000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel126[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel126_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel126 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111101000011000110001001001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel126[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel126_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel126 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111110000010111001111101010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel126[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel126_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel126 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b10111100100001001000100101011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel126[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel126_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel126 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b10111110101010001110010101011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel126[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel126_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel126 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111110100011001110111101001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel126[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel126_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel126 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b00111100111010101110001101101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel126[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel126_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel126 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b10111100111101001110000111010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel126[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel126_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel126 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b10111100101110010000001011011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel126[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel126_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel126 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b10111110001111011011010111001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel126[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel126_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel126 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b10111110101100100001100000111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel126[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel126_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel126 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111100010010100010001101001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel126[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel126_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel126 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111101010011011100111110100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel126[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel126_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel126 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b10111100001011110000010011000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel126[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel126_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel126 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111101011010001110010001100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel126[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel126_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel126 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b10111110100010010000000000011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel126[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel126_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel126 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111110100110110001101110100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel126[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel126_Valid_Out)
	);
	Adder_64input add_k126(
		.Data1(Data_Out_Kernel126[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel126[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel126[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel126[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel126[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel126[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel126[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel126[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel126[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel126[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel126[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel126[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel126[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel126[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel126[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel126[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel126[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel126[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel126[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel126[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel126[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel126[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel126[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel126[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel126[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel126[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel126[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel126[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel126[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel126[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel126[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel126[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel126[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel126[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel126[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel126[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel126[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel126[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel126[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel126[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel126[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel126[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel126[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel126[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel126[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel126[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel126[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel126[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel126[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel126[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel126[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel126[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel126[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel126[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel126[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel126[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel126[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel126[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel126[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel126[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel126[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel126[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel126[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel126[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel126),
		.Data_Out(add_k126_Data_Out),
		.Valid_Out(add_kernel126_Valid_Out)
	);
	Batch_Norm bn_kernel126(
		.Data_A(32'b00111110010110011100101010101011),
		.Data_B(32'b00111110101010111010110000101001),
		.Data_In(add_k126_Data_Out),
		.Valid_In(add_kernel126_Valid_Out),
		.Data_Out(bn126_Data_Out),
		.Valid_Out(bn126_Valid_Out)
	);
	Relu_Core rl_kernel126(
		.Data_In(bn126_Data_Out),
		.Valid_In(bn126_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*126-1:DATA_WIDHT*125]),
		.Valid_Out(rl126_Valid_Out)
	);
//////////KERNEL127//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel127 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111111000000010011111100100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel127[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel127_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel127 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110001101101010011111110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel127[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel127_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel127 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111101011101100101011001110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel127[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel127_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel127 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111111000010101010000111101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel127[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel127_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel127 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111101100110011110011101101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel127[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel127_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel127 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110010001000011100111110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel127[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel127_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel127 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111101101010001011110100100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel127[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel127_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel127 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111101100000100011011001010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel127[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel127_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel127 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111101001101111110101110111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel127[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel127_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel127 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111101110001011100001001110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel127[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel127_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel127 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111101101000010110110011011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel127[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel127_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel127 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111101111000001000001011100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel127[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel127_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel127 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110000010100111100110100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel127[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel127_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel127 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111100111011101001110001001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel127[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel127_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel127 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111101101011001010001100001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel127[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel127_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel127 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111100111111111111111100100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel127[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel127_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel127 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111101010000000101110110011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel127[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel127_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel127 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111101111110100011110100101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel127[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel127_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel127 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110011010010101001011100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel127[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel127_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel127 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111101110111100101110101110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel127[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel127_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel127 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111111000000111010000111111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel127[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel127_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel127 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111110001001111111110010100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel127[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel127_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel127 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111111001010000011000000001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel127[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel127_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel127 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111111000000000100000111110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel127[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel127_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel127 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111110111001101001111010101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel127[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel127_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel127 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110110101101001100110101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel127[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel127_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel127 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110100010001010111011101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel127[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel127_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel127 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111110000100011111110001000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel127[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel127_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel127 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111110111010010111110100110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel127[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel127_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel127 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111110101011100110000101110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel127[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel127_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel127 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111101110010100110100111101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel127[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel127_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel127 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110111111010101100001110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel127[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel127_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel127 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111110101100100100010000000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel127[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel127_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel127 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b10111101100100101100101101101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel127[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel127_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel127 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111110011110111011110101001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel127[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel127_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel127 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111110010011001101011001110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel127[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel127_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel127 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111110101111111011111001101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel127[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel127_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel127 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b00111101110000010001101111101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel127[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel127_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel127 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b00111111000110001011110000000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel127[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel127_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel127 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111110100011111011110100101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel127[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel127_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel127 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111111010001111101000110100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel127[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel127_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel127 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111110100101010001110100110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel127[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel127_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel127 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b10111110101101000001111010010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel127[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel127_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel127 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b00111110111100110011110101000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel127[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel127_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel127 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111111000101001111001001001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel127[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel127_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel127 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111110010011111010011110111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel127[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel127_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel127 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b10111110011011111100011001110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel127[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel127_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel127 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111101000011000000011110111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel127[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel127_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel127 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111110101011010000100110011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel127[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel127_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel127 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b10111101100101111110111110010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel127[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel127_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel127 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111110110111110100011010011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel127[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel127_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel127 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111110011011101101000101000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel127[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel127_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel127 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b10111110010111101001101101011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel127[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel127_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel127 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111111000111101100111000100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel127[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel127_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel127 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b00111110011111011011001001100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel127[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel127_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel127 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b00111100001001001000010011100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel127[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel127_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel127 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111101011101111010110110010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel127[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel127_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel127 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b00111110011001111110111100011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel127[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel127_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel127 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b00111110000110101100001101110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel127[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel127_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel127 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111110111000111011011010010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel127[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel127_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel127 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111110101111100101001110110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel127[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel127_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel127 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111101100101101101000001101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel127[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel127_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel127 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111111000101010000110100001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel127[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel127_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel127 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b10111110110011110001110000001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel127[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel127_Valid_Out)
	);
	Adder_64input add_k127(
		.Data1(Data_Out_Kernel127[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel127[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel127[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel127[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel127[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel127[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel127[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel127[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel127[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel127[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel127[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel127[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel127[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel127[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel127[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel127[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel127[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel127[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel127[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel127[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel127[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel127[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel127[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel127[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel127[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel127[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel127[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel127[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel127[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel127[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel127[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel127[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel127[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel127[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel127[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel127[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel127[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel127[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel127[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel127[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel127[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel127[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel127[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel127[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel127[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel127[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel127[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel127[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel127[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel127[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel127[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel127[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel127[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel127[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel127[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel127[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel127[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel127[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel127[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel127[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel127[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel127[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel127[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel127[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel127),
		.Data_Out(add_k127_Data_Out),
		.Valid_Out(add_kernel127_Valid_Out)
	);
	Batch_Norm bn_kernel127(
		.Data_A(32'b00111110000100001100000100100111),
		.Data_B(32'b10111110110011001011001010111000),
		.Data_In(add_k127_Data_Out),
		.Valid_In(add_kernel127_Valid_Out),
		.Data_Out(bn127_Data_Out),
		.Valid_Out(bn127_Valid_Out)
	);
	Relu_Core rl_kernel127(
		.Data_In(bn127_Data_Out),
		.Valid_In(bn127_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*127-1:DATA_WIDHT*126]),
		.Valid_Out(rl127_Valid_Out)
	);
//////////KERNEL128//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel128 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111110111110001010010011011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel128[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel128_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel128 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111101111111011001010100000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel128[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel128_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel128 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110000101100001111000011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel128[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel128_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel128 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110100111011111101101111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel128[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel128_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel128 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111110010100000110100111000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel128[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel128_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel128 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111101011101011011110101010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel128[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel128_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel128 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111101100110110110101101011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel128[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel128_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel128 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111101100110100000101111101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel128[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel128_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel128 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111100110001101001111101111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel128[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel128_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel128 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111100100110111000001000000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel128[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel128_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel128 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111100111001100010110010100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel128[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel128_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel128 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111110001001011000110001100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel128[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel128_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel128 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110000000110011111111010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel128[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel128_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel128 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111110001111100000011011101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel128[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel128_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel128 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110110000010111000011001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel128[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel128_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel128 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111101000011101010000100101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel128[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel128_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel128 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111111000110111001100011010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel128[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel128_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel128 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111101001011000011010010111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel128[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel128_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel128 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111101100111000011110111001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel128[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel128_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel128 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110001011000100010101001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel128[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel128_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel128 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110100000000001110110111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel128[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel128_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel128 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111101111001110111010011011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel128[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel128_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel128 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111101111101100101111100001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel128[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel128_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel128 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111110010011001010001111001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel128[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel128_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel128 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111110101111111011001000001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel128[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel128_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel128 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110100100101011101011000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel128[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel128_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel128 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110010100111001100101010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel128[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel128_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel128 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111110010000111010111000011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel128[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel128_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel128 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111110010101010101110101101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel128[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel128_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel128 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111100000000000010011000101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel128[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel128_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel128 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111110001000010001010100111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel128[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel128_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel128 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110101110101011100110101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel128[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel128_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL33_Kernel128 (
		.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Kernel(32'b10111110000001011000000101110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel128[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(channel33_Kernel128_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL34_Kernel128 (
		.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Kernel(32'b00111101001010010110100111011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel128[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(channel34_Kernel128_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL35_Kernel128 (
		.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Kernel(32'b00111110101000000100100111110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel128[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(channel35_Kernel128_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL36_Kernel128 (
		.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Kernel(32'b00111100000110000110000010110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel128[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(channel36_Kernel128_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL37_Kernel128 (
		.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Kernel(32'b00111110011110010001000010110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel128[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(channel37_Kernel128_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL38_Kernel128 (
		.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Kernel(32'b00111100110010010111001011010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel128[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(channel38_Kernel128_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL39_Kernel128 (
		.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Kernel(32'b00111110011001011000110000011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel128[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(channel39_Kernel128_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL40_Kernel128 (
		.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Kernel(32'b10111110001000100100001000000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel128[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(channel40_Kernel128_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL41_Kernel128 (
		.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Kernel(32'b00111111000111000000001000000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel128[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(channel41_Kernel128_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL42_Kernel128 (
		.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Kernel(32'b00111110101100010011101011100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel128[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(channel42_Kernel128_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL43_Kernel128 (
		.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Kernel(32'b00111010101100000111101111010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel128[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(channel43_Kernel128_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL44_Kernel128 (
		.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Kernel(32'b00111100011101010010100010010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel128[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(channel44_Kernel128_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL45_Kernel128 (
		.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Kernel(32'b10111110100010110010101110110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel128[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(channel45_Kernel128_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL46_Kernel128 (
		.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Kernel(32'b00111110001110000100010011010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel128[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(channel46_Kernel128_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL47_Kernel128 (
		.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Kernel(32'b00111110011101111110001000101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel128[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(channel47_Kernel128_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL48_Kernel128 (
		.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Kernel(32'b10111110100001110111110101001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel128[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(channel48_Kernel128_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL49_Kernel128 (
		.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Kernel(32'b10111101110010000101010110110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel128[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(channel49_Kernel128_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL50_Kernel128 (
		.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Kernel(32'b00111100001100111001100110011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel128[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(channel50_Kernel128_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL51_Kernel128 (
		.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Kernel(32'b00111110011110110101001000000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel128[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(channel51_Kernel128_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL52_Kernel128 (
		.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Kernel(32'b00111101010011110001110110010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel128[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(channel52_Kernel128_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL53_Kernel128 (
		.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Kernel(32'b00111110001011100010110100101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel128[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(channel53_Kernel128_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL54_Kernel128 (
		.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Kernel(32'b10111110111110011001100111100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel128[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(channel54_Kernel128_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL55_Kernel128 (
		.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Kernel(32'b10111110000000011100100000100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel128[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(channel55_Kernel128_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL56_Kernel128 (
		.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Kernel(32'b00111011001011100110000101110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel128[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(channel56_Kernel128_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL57_Kernel128 (
		.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Kernel(32'b00111110110010001101000101110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel128[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(channel57_Kernel128_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL58_Kernel128 (
		.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Kernel(32'b10111100100011100011100011011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel128[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(channel58_Kernel128_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL59_Kernel128 (
		.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Kernel(32'b10111100101100010111100010111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel128[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(channel59_Kernel128_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL60_Kernel128 (
		.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Kernel(32'b10111011100110001101110101100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel128[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(channel60_Kernel128_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL61_Kernel128 (
		.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Kernel(32'b00111110001101011001110110110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel128[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(channel61_Kernel128_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL62_Kernel128 (
		.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Kernel(32'b00111101010110110100001100000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel128[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(channel62_Kernel128_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL63_Kernel128 (
		.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Kernel(32'b00111101101110110100001010001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel128[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(channel63_Kernel128_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL64_Kernel128 (
		.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Kernel(32'b00111011100101001110010010011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel128[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(channel64_Kernel128_Valid_Out)
	);
	Adder_64input add_k128(
		.Data1(Data_Out_Kernel128[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel128[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel128[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel128[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel128[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel128[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel128[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel128[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel128[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel128[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel128[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel128[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel128[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel128[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel128[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel128[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel128[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel128[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel128[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel128[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel128[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel128[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel128[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel128[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel128[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel128[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel128[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel128[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel128[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel128[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel128[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel128[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Data33(Data_Out_Kernel128[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Data34(Data_Out_Kernel128[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Data35(Data_Out_Kernel128[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Data36(Data_Out_Kernel128[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Data37(Data_Out_Kernel128[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Data38(Data_Out_Kernel128[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Data39(Data_Out_Kernel128[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Data40(Data_Out_Kernel128[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Data41(Data_Out_Kernel128[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Data42(Data_Out_Kernel128[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Data43(Data_Out_Kernel128[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Data44(Data_Out_Kernel128[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Data45(Data_Out_Kernel128[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Data46(Data_Out_Kernel128[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Data47(Data_Out_Kernel128[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Data48(Data_Out_Kernel128[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Data49(Data_Out_Kernel128[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Data50(Data_Out_Kernel128[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Data51(Data_Out_Kernel128[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Data52(Data_Out_Kernel128[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Data53(Data_Out_Kernel128[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Data54(Data_Out_Kernel128[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Data55(Data_Out_Kernel128[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Data56(Data_Out_Kernel128[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Data57(Data_Out_Kernel128[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Data58(Data_Out_Kernel128[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Data59(Data_Out_Kernel128[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Data60(Data_Out_Kernel128[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Data61(Data_Out_Kernel128[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Data62(Data_Out_Kernel128[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Data63(Data_Out_Kernel128[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Data64(Data_Out_Kernel128[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_In(add_kernel128),
		.Data_Out(add_k128_Data_Out),
		.Valid_Out(add_kernel128_Valid_Out)
	);
	Batch_Norm bn_kernel128(
		.Data_A(32'b00111110010011000010001001011001),
		.Data_B(32'b10111111010000110101011001000000),
		.Data_In(add_k128_Data_Out),
		.Valid_In(add_kernel128_Valid_Out),
		.Data_Out(bn128_Data_Out),
		.Valid_Out(bn128_Valid_Out)
	);
	Relu_Core rl_kernel128(
		.Data_In(bn128_Data_Out),
		.Valid_In(bn128_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*128-1:DATA_WIDHT*127]),
		.Valid_Out(rl128_Valid_Out)
	);

    
endmodule