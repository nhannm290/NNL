module Layer6 #(
    parameter DATA_WIDHT = 32,
    parameter IMG_WIDHT = 44,
    parameter IMG_HEIGHT =44
)

(
    input [DATA_WIDHT*64-1:0] Data_In,
    input clk,
    input rst,
    input Valid_In,
    output [DATA_WIDHT*128-1:0] Data_Out,
    output Valid_Out    
);

    wire [DATA_WIDHT*128-1:0] sp_8Channel_Data_Out,sp_16Channel_Data_Out,Convo3_Data_Out,lb_Data_Out,Max_Data_Out;
    wire sp_8Channel_Valid_Out,sp_16Channel_Valid_Out,Convo_Valid_Out,lb_Valid_Out,add_Valid_In,Max_Valid_Out;

    assign add_Valid_In = Max_Valid_Out& lb_Valid_Out;


    Separable_Convolution_Part1_Layer6 #(
        .DATA_WIDHT(DATA_WIDHT),
        .IMG_WIDHT(IMG_WIDHT),
        .IMG_HEIGHT(IMG_HEIGHT)
    )
        sp_convo_16channel (
            .Data_In(Data_In),
            .Valid_In(Valid_In),
            .clk(clk),
            .rst(rst),
            .Data_Out(sp_8Channel_Data_Out),
            .Valid_Out(sp_8Channel_Valid_Out)
        );

    Separable_Convolution_Part2_Layer6 #(
        .DATA_WIDHT(DATA_WIDHT),
        .IMG_WIDHT(IMG_WIDHT),
        .IMG_HEIGHT(IMG_HEIGHT)
    )
        sp_convo_32channel(
            .Data_In(sp_8Channel_Data_Out),
            .Valid_In(sp_8Channel_Valid_Out),
            .clk(clk),
            .rst(rst),
            .Data_Out(sp_16Channel_Data_Out),
            .Valid_Out(sp_16Channel_Valid_Out)
        );

    MaxPooling_3x3_stride_1x1_padding_1 #(
        .DATA_WIDHT(DATA_WIDHT),
        .IMG_WIDHT(IMG_WIDHT),
        .IMG_HEIGHT(IMG_HEIGHT)
    )   
        maxpooling[127:0] (
            .Data_In({sp_16Channel_Data_Out[DATA_WIDHT-1:0], sp_16Channel_Data_Out[DATA_WIDHT*2-1:DATA_WIDHT],sp_16Channel_Data_Out[DATA_WIDHT*3-1:DATA_WIDHT*2],sp_16Channel_Data_Out[DATA_WIDHT*4-1:DATA_WIDHT*3],sp_16Channel_Data_Out[DATA_WIDHT*5-1:DATA_WIDHT*4],sp_16Channel_Data_Out[DATA_WIDHT*6-1:DATA_WIDHT*5],sp_16Channel_Data_Out[DATA_WIDHT*7-1:DATA_WIDHT*6],sp_16Channel_Data_Out[DATA_WIDHT*8-1:DATA_WIDHT*7],sp_16Channel_Data_Out[DATA_WIDHT*9-1:DATA_WIDHT*8],sp_16Channel_Data_Out[DATA_WIDHT*10-1:DATA_WIDHT*9],sp_16Channel_Data_Out[DATA_WIDHT*11-1:DATA_WIDHT*10],sp_16Channel_Data_Out[DATA_WIDHT*12-1:DATA_WIDHT*11],sp_16Channel_Data_Out[DATA_WIDHT*13-1:DATA_WIDHT*12],sp_16Channel_Data_Out[DATA_WIDHT*14-1:DATA_WIDHT*13],sp_16Channel_Data_Out[DATA_WIDHT*15-1:DATA_WIDHT*14],sp_16Channel_Data_Out[DATA_WIDHT*16-1:DATA_WIDHT*15],sp_16Channel_Data_Out[DATA_WIDHT*17-1:DATA_WIDHT*16],sp_16Channel_Data_Out[DATA_WIDHT*18-1:DATA_WIDHT*17],sp_16Channel_Data_Out[DATA_WIDHT*19-1:DATA_WIDHT*18],sp_16Channel_Data_Out[DATA_WIDHT*20-1:DATA_WIDHT*19],sp_16Channel_Data_Out[DATA_WIDHT*21-1:DATA_WIDHT*20],sp_16Channel_Data_Out[DATA_WIDHT*22-1:DATA_WIDHT*21],sp_16Channel_Data_Out[DATA_WIDHT*23-1:DATA_WIDHT*22],sp_16Channel_Data_Out[DATA_WIDHT*24-1:DATA_WIDHT*23],sp_16Channel_Data_Out[DATA_WIDHT*25-1:DATA_WIDHT*24],sp_16Channel_Data_Out[DATA_WIDHT*26-1:DATA_WIDHT*25],sp_16Channel_Data_Out[DATA_WIDHT*27-1:DATA_WIDHT*26],sp_16Channel_Data_Out[DATA_WIDHT*28-1:DATA_WIDHT*27],sp_16Channel_Data_Out[DATA_WIDHT*29-1:DATA_WIDHT*28],sp_16Channel_Data_Out[DATA_WIDHT*30-1:DATA_WIDHT*29],sp_16Channel_Data_Out[DATA_WIDHT*31-1:DATA_WIDHT*30],sp_16Channel_Data_Out[DATA_WIDHT*32-1:DATA_WIDHT*31],sp_16Channel_Data_Out[DATA_WIDHT*33-1:DATA_WIDHT*32],sp_16Channel_Data_Out[DATA_WIDHT*34-1:DATA_WIDHT*33],sp_16Channel_Data_Out[DATA_WIDHT*35-1:DATA_WIDHT*34],sp_16Channel_Data_Out[DATA_WIDHT*36-1:DATA_WIDHT*35],sp_16Channel_Data_Out[DATA_WIDHT*37-1:DATA_WIDHT*36],sp_16Channel_Data_Out[DATA_WIDHT*38-1:DATA_WIDHT*37],sp_16Channel_Data_Out[DATA_WIDHT*39-1:DATA_WIDHT*38],sp_16Channel_Data_Out[DATA_WIDHT*40-1:DATA_WIDHT*39],sp_16Channel_Data_Out[DATA_WIDHT*41-1:DATA_WIDHT*40],sp_16Channel_Data_Out[DATA_WIDHT*42-1:DATA_WIDHT*41],sp_16Channel_Data_Out[DATA_WIDHT*43-1:DATA_WIDHT*42],sp_16Channel_Data_Out[DATA_WIDHT*44-1:DATA_WIDHT*43],sp_16Channel_Data_Out[DATA_WIDHT*45-1:DATA_WIDHT*44],sp_16Channel_Data_Out[DATA_WIDHT*46-1:DATA_WIDHT*45],sp_16Channel_Data_Out[DATA_WIDHT*47-1:DATA_WIDHT*46],sp_16Channel_Data_Out[DATA_WIDHT*48-1:DATA_WIDHT*47],sp_16Channel_Data_Out[DATA_WIDHT*49-1:DATA_WIDHT*48],sp_16Channel_Data_Out[DATA_WIDHT*50-1:DATA_WIDHT*49],sp_16Channel_Data_Out[DATA_WIDHT*51-1:DATA_WIDHT*50],sp_16Channel_Data_Out[DATA_WIDHT*52-1:DATA_WIDHT*51],sp_16Channel_Data_Out[DATA_WIDHT*53-1:DATA_WIDHT*52],sp_16Channel_Data_Out[DATA_WIDHT*54-1:DATA_WIDHT*53],sp_16Channel_Data_Out[DATA_WIDHT*55-1:DATA_WIDHT*54],sp_16Channel_Data_Out[DATA_WIDHT*56-1:DATA_WIDHT*55],sp_16Channel_Data_Out[DATA_WIDHT*57-1:DATA_WIDHT*56],sp_16Channel_Data_Out[DATA_WIDHT*58-1:DATA_WIDHT*57],sp_16Channel_Data_Out[DATA_WIDHT*59-1:DATA_WIDHT*58],sp_16Channel_Data_Out[DATA_WIDHT*60-1:DATA_WIDHT*59],sp_16Channel_Data_Out[DATA_WIDHT*61-1:DATA_WIDHT*60],sp_16Channel_Data_Out[DATA_WIDHT*62-1:DATA_WIDHT*61],sp_16Channel_Data_Out[DATA_WIDHT*63-1:DATA_WIDHT*62],sp_16Channel_Data_Out[DATA_WIDHT*64-1:DATA_WIDHT*63],sp_16Channel_Data_Out[DATA_WIDHT*65-1:DATA_WIDHT*64],sp_16Channel_Data_Out[DATA_WIDHT*66-1:DATA_WIDHT*65],sp_16Channel_Data_Out[DATA_WIDHT*67-1:DATA_WIDHT*66],sp_16Channel_Data_Out[DATA_WIDHT*68-1:DATA_WIDHT*67],sp_16Channel_Data_Out[DATA_WIDHT*69-1:DATA_WIDHT*68],sp_16Channel_Data_Out[DATA_WIDHT*70-1:DATA_WIDHT*69],sp_16Channel_Data_Out[DATA_WIDHT*71-1:DATA_WIDHT*70],sp_16Channel_Data_Out[DATA_WIDHT*72-1:DATA_WIDHT*71],sp_16Channel_Data_Out[DATA_WIDHT*73-1:DATA_WIDHT*72],sp_16Channel_Data_Out[DATA_WIDHT*74-1:DATA_WIDHT*73],sp_16Channel_Data_Out[DATA_WIDHT*75-1:DATA_WIDHT*74],sp_16Channel_Data_Out[DATA_WIDHT*76-1:DATA_WIDHT*75],sp_16Channel_Data_Out[DATA_WIDHT*77-1:DATA_WIDHT*76],sp_16Channel_Data_Out[DATA_WIDHT*78-1:DATA_WIDHT*77],sp_16Channel_Data_Out[DATA_WIDHT*79-1:DATA_WIDHT*78],sp_16Channel_Data_Out[DATA_WIDHT*80-1:DATA_WIDHT*79],sp_16Channel_Data_Out[DATA_WIDHT*81-1:DATA_WIDHT*80],sp_16Channel_Data_Out[DATA_WIDHT*82-1:DATA_WIDHT*81],sp_16Channel_Data_Out[DATA_WIDHT*83-1:DATA_WIDHT*82],sp_16Channel_Data_Out[DATA_WIDHT*84-1:DATA_WIDHT*83],sp_16Channel_Data_Out[DATA_WIDHT*85-1:DATA_WIDHT*84],sp_16Channel_Data_Out[DATA_WIDHT*86-1:DATA_WIDHT*85],sp_16Channel_Data_Out[DATA_WIDHT*87-1:DATA_WIDHT*86],sp_16Channel_Data_Out[DATA_WIDHT*88-1:DATA_WIDHT*87],sp_16Channel_Data_Out[DATA_WIDHT*89-1:DATA_WIDHT*88],sp_16Channel_Data_Out[DATA_WIDHT*90-1:DATA_WIDHT*89],sp_16Channel_Data_Out[DATA_WIDHT*91-1:DATA_WIDHT*90],sp_16Channel_Data_Out[DATA_WIDHT*92-1:DATA_WIDHT*91],sp_16Channel_Data_Out[DATA_WIDHT*93-1:DATA_WIDHT*92],sp_16Channel_Data_Out[DATA_WIDHT*94-1:DATA_WIDHT*93],sp_16Channel_Data_Out[DATA_WIDHT*95-1:DATA_WIDHT*94],sp_16Channel_Data_Out[DATA_WIDHT*96-1:DATA_WIDHT*95],sp_16Channel_Data_Out[DATA_WIDHT*97-1:DATA_WIDHT*96],sp_16Channel_Data_Out[DATA_WIDHT*98-1:DATA_WIDHT*97],sp_16Channel_Data_Out[DATA_WIDHT*99-1:DATA_WIDHT*98],sp_16Channel_Data_Out[DATA_WIDHT*100-1:DATA_WIDHT*99],sp_16Channel_Data_Out[DATA_WIDHT*101-1:DATA_WIDHT*100],sp_16Channel_Data_Out[DATA_WIDHT*102-1:DATA_WIDHT*101],sp_16Channel_Data_Out[DATA_WIDHT*103-1:DATA_WIDHT*102],sp_16Channel_Data_Out[DATA_WIDHT*104-1:DATA_WIDHT*103],sp_16Channel_Data_Out[DATA_WIDHT*105-1:DATA_WIDHT*104],sp_16Channel_Data_Out[DATA_WIDHT*106-1:DATA_WIDHT*105],sp_16Channel_Data_Out[DATA_WIDHT*107-1:DATA_WIDHT*106],sp_16Channel_Data_Out[DATA_WIDHT*108-1:DATA_WIDHT*107],sp_16Channel_Data_Out[DATA_WIDHT*109-1:DATA_WIDHT*108],sp_16Channel_Data_Out[DATA_WIDHT*110-1:DATA_WIDHT*109],sp_16Channel_Data_Out[DATA_WIDHT*111-1:DATA_WIDHT*110],sp_16Channel_Data_Out[DATA_WIDHT*112-1:DATA_WIDHT*111],sp_16Channel_Data_Out[DATA_WIDHT*113-1:DATA_WIDHT*112],sp_16Channel_Data_Out[DATA_WIDHT*114-1:DATA_WIDHT*113],sp_16Channel_Data_Out[DATA_WIDHT*115-1:DATA_WIDHT*114],sp_16Channel_Data_Out[DATA_WIDHT*116-1:DATA_WIDHT*115],sp_16Channel_Data_Out[DATA_WIDHT*117-1:DATA_WIDHT*116],sp_16Channel_Data_Out[DATA_WIDHT*118-1:DATA_WIDHT*117],sp_16Channel_Data_Out[DATA_WIDHT*119-1:DATA_WIDHT*118],sp_16Channel_Data_Out[DATA_WIDHT*120-1:DATA_WIDHT*119],sp_16Channel_Data_Out[DATA_WIDHT*121-1:DATA_WIDHT*120],sp_16Channel_Data_Out[DATA_WIDHT*122-1:DATA_WIDHT*121],sp_16Channel_Data_Out[DATA_WIDHT*123-1:DATA_WIDHT*122],sp_16Channel_Data_Out[DATA_WIDHT*124-1:DATA_WIDHT*123],sp_16Channel_Data_Out[DATA_WIDHT*125-1:DATA_WIDHT*124],sp_16Channel_Data_Out[DATA_WIDHT*126-1:DATA_WIDHT*125],sp_16Channel_Data_Out[DATA_WIDHT*127-1:DATA_WIDHT*126],sp_16Channel_Data_Out[DATA_WIDHT*128-1:DATA_WIDHT*127]}),
            .Valid_In(sp_16Channel_Valid_Out),
            .clk(clk),
            .rst(rst),
            .Data_Out({Max_Data_Out[DATA_WIDHT-1:0], Max_Data_Out[DATA_WIDHT*2-1:DATA_WIDHT],Max_Data_Out[DATA_WIDHT*3-1:DATA_WIDHT*2],Max_Data_Out[DATA_WIDHT*4-1:DATA_WIDHT*3],Max_Data_Out[DATA_WIDHT*5-1:DATA_WIDHT*4],Max_Data_Out[DATA_WIDHT*6-1:DATA_WIDHT*5],Max_Data_Out[DATA_WIDHT*7-1:DATA_WIDHT*6],Max_Data_Out[DATA_WIDHT*8-1:DATA_WIDHT*7],Max_Data_Out[DATA_WIDHT*9-1:DATA_WIDHT*8],Max_Data_Out[DATA_WIDHT*10-1:DATA_WIDHT*9],Max_Data_Out[DATA_WIDHT*11-1:DATA_WIDHT*10],Max_Data_Out[DATA_WIDHT*12-1:DATA_WIDHT*11],Max_Data_Out[DATA_WIDHT*13-1:DATA_WIDHT*12],Max_Data_Out[DATA_WIDHT*14-1:DATA_WIDHT*13],Max_Data_Out[DATA_WIDHT*15-1:DATA_WIDHT*14],Max_Data_Out[DATA_WIDHT*16-1:DATA_WIDHT*15],Max_Data_Out[DATA_WIDHT*17-1:DATA_WIDHT*16],Max_Data_Out[DATA_WIDHT*18-1:DATA_WIDHT*17],Max_Data_Out[DATA_WIDHT*19-1:DATA_WIDHT*18],Max_Data_Out[DATA_WIDHT*20-1:DATA_WIDHT*19],Max_Data_Out[DATA_WIDHT*21-1:DATA_WIDHT*20],Max_Data_Out[DATA_WIDHT*22-1:DATA_WIDHT*21],Max_Data_Out[DATA_WIDHT*23-1:DATA_WIDHT*22],Max_Data_Out[DATA_WIDHT*24-1:DATA_WIDHT*23],Max_Data_Out[DATA_WIDHT*25-1:DATA_WIDHT*24],Max_Data_Out[DATA_WIDHT*26-1:DATA_WIDHT*25],Max_Data_Out[DATA_WIDHT*27-1:DATA_WIDHT*26],Max_Data_Out[DATA_WIDHT*28-1:DATA_WIDHT*27],Max_Data_Out[DATA_WIDHT*29-1:DATA_WIDHT*28],Max_Data_Out[DATA_WIDHT*30-1:DATA_WIDHT*29],Max_Data_Out[DATA_WIDHT*31-1:DATA_WIDHT*30],Max_Data_Out[DATA_WIDHT*32-1:DATA_WIDHT*31],Max_Data_Out[DATA_WIDHT*33-1:DATA_WIDHT*32],Max_Data_Out[DATA_WIDHT*34-1:DATA_WIDHT*33],Max_Data_Out[DATA_WIDHT*35-1:DATA_WIDHT*34],Max_Data_Out[DATA_WIDHT*36-1:DATA_WIDHT*35],Max_Data_Out[DATA_WIDHT*37-1:DATA_WIDHT*36],Max_Data_Out[DATA_WIDHT*38-1:DATA_WIDHT*37],Max_Data_Out[DATA_WIDHT*39-1:DATA_WIDHT*38],Max_Data_Out[DATA_WIDHT*40-1:DATA_WIDHT*39],Max_Data_Out[DATA_WIDHT*41-1:DATA_WIDHT*40],Max_Data_Out[DATA_WIDHT*42-1:DATA_WIDHT*41],Max_Data_Out[DATA_WIDHT*43-1:DATA_WIDHT*42],Max_Data_Out[DATA_WIDHT*44-1:DATA_WIDHT*43],Max_Data_Out[DATA_WIDHT*45-1:DATA_WIDHT*44],Max_Data_Out[DATA_WIDHT*46-1:DATA_WIDHT*45],Max_Data_Out[DATA_WIDHT*47-1:DATA_WIDHT*46],Max_Data_Out[DATA_WIDHT*48-1:DATA_WIDHT*47],Max_Data_Out[DATA_WIDHT*49-1:DATA_WIDHT*48],Max_Data_Out[DATA_WIDHT*50-1:DATA_WIDHT*49],Max_Data_Out[DATA_WIDHT*51-1:DATA_WIDHT*50],Max_Data_Out[DATA_WIDHT*52-1:DATA_WIDHT*51],Max_Data_Out[DATA_WIDHT*53-1:DATA_WIDHT*52],Max_Data_Out[DATA_WIDHT*54-1:DATA_WIDHT*53],Max_Data_Out[DATA_WIDHT*55-1:DATA_WIDHT*54],Max_Data_Out[DATA_WIDHT*56-1:DATA_WIDHT*55],Max_Data_Out[DATA_WIDHT*57-1:DATA_WIDHT*56],Max_Data_Out[DATA_WIDHT*58-1:DATA_WIDHT*57],Max_Data_Out[DATA_WIDHT*59-1:DATA_WIDHT*58],Max_Data_Out[DATA_WIDHT*60-1:DATA_WIDHT*59],Max_Data_Out[DATA_WIDHT*61-1:DATA_WIDHT*60],Max_Data_Out[DATA_WIDHT*62-1:DATA_WIDHT*61],Max_Data_Out[DATA_WIDHT*63-1:DATA_WIDHT*62],Max_Data_Out[DATA_WIDHT*64-1:DATA_WIDHT*63],Max_Data_Out[DATA_WIDHT*65-1:DATA_WIDHT*64],Max_Data_Out[DATA_WIDHT*66-1:DATA_WIDHT*65],Max_Data_Out[DATA_WIDHT*67-1:DATA_WIDHT*66],Max_Data_Out[DATA_WIDHT*68-1:DATA_WIDHT*67],Max_Data_Out[DATA_WIDHT*69-1:DATA_WIDHT*68],Max_Data_Out[DATA_WIDHT*70-1:DATA_WIDHT*69],Max_Data_Out[DATA_WIDHT*71-1:DATA_WIDHT*70],Max_Data_Out[DATA_WIDHT*72-1:DATA_WIDHT*71],Max_Data_Out[DATA_WIDHT*73-1:DATA_WIDHT*72],Max_Data_Out[DATA_WIDHT*74-1:DATA_WIDHT*73],Max_Data_Out[DATA_WIDHT*75-1:DATA_WIDHT*74],Max_Data_Out[DATA_WIDHT*76-1:DATA_WIDHT*75],Max_Data_Out[DATA_WIDHT*77-1:DATA_WIDHT*76],Max_Data_Out[DATA_WIDHT*78-1:DATA_WIDHT*77],Max_Data_Out[DATA_WIDHT*79-1:DATA_WIDHT*78],Max_Data_Out[DATA_WIDHT*80-1:DATA_WIDHT*79],Max_Data_Out[DATA_WIDHT*81-1:DATA_WIDHT*80],Max_Data_Out[DATA_WIDHT*82-1:DATA_WIDHT*81],Max_Data_Out[DATA_WIDHT*83-1:DATA_WIDHT*82],Max_Data_Out[DATA_WIDHT*84-1:DATA_WIDHT*83],Max_Data_Out[DATA_WIDHT*85-1:DATA_WIDHT*84],Max_Data_Out[DATA_WIDHT*86-1:DATA_WIDHT*85],Max_Data_Out[DATA_WIDHT*87-1:DATA_WIDHT*86],Max_Data_Out[DATA_WIDHT*88-1:DATA_WIDHT*87],Max_Data_Out[DATA_WIDHT*89-1:DATA_WIDHT*88],Max_Data_Out[DATA_WIDHT*90-1:DATA_WIDHT*89],Max_Data_Out[DATA_WIDHT*91-1:DATA_WIDHT*90],Max_Data_Out[DATA_WIDHT*92-1:DATA_WIDHT*91],Max_Data_Out[DATA_WIDHT*93-1:DATA_WIDHT*92],Max_Data_Out[DATA_WIDHT*94-1:DATA_WIDHT*93],Max_Data_Out[DATA_WIDHT*95-1:DATA_WIDHT*94],Max_Data_Out[DATA_WIDHT*96-1:DATA_WIDHT*95],Max_Data_Out[DATA_WIDHT*97-1:DATA_WIDHT*96],Max_Data_Out[DATA_WIDHT*98-1:DATA_WIDHT*97],Max_Data_Out[DATA_WIDHT*99-1:DATA_WIDHT*98],Max_Data_Out[DATA_WIDHT*100-1:DATA_WIDHT*99],Max_Data_Out[DATA_WIDHT*101-1:DATA_WIDHT*100],Max_Data_Out[DATA_WIDHT*102-1:DATA_WIDHT*101],Max_Data_Out[DATA_WIDHT*103-1:DATA_WIDHT*102],Max_Data_Out[DATA_WIDHT*104-1:DATA_WIDHT*103],Max_Data_Out[DATA_WIDHT*105-1:DATA_WIDHT*104],Max_Data_Out[DATA_WIDHT*106-1:DATA_WIDHT*105],Max_Data_Out[DATA_WIDHT*107-1:DATA_WIDHT*106],Max_Data_Out[DATA_WIDHT*108-1:DATA_WIDHT*107],Max_Data_Out[DATA_WIDHT*109-1:DATA_WIDHT*108],Max_Data_Out[DATA_WIDHT*110-1:DATA_WIDHT*109],Max_Data_Out[DATA_WIDHT*111-1:DATA_WIDHT*110],Max_Data_Out[DATA_WIDHT*112-1:DATA_WIDHT*111],Max_Data_Out[DATA_WIDHT*113-1:DATA_WIDHT*112],Max_Data_Out[DATA_WIDHT*114-1:DATA_WIDHT*113],Max_Data_Out[DATA_WIDHT*115-1:DATA_WIDHT*114],Max_Data_Out[DATA_WIDHT*116-1:DATA_WIDHT*115],Max_Data_Out[DATA_WIDHT*117-1:DATA_WIDHT*116],Max_Data_Out[DATA_WIDHT*118-1:DATA_WIDHT*117],Max_Data_Out[DATA_WIDHT*119-1:DATA_WIDHT*118],Max_Data_Out[DATA_WIDHT*120-1:DATA_WIDHT*119],Max_Data_Out[DATA_WIDHT*121-1:DATA_WIDHT*120],Max_Data_Out[DATA_WIDHT*122-1:DATA_WIDHT*121],Max_Data_Out[DATA_WIDHT*123-1:DATA_WIDHT*122],Max_Data_Out[DATA_WIDHT*124-1:DATA_WIDHT*123],Max_Data_Out[DATA_WIDHT*125-1:DATA_WIDHT*124],Max_Data_Out[DATA_WIDHT*126-1:DATA_WIDHT*125],Max_Data_Out[DATA_WIDHT*127-1:DATA_WIDHT*126],Max_Data_Out[DATA_WIDHT*128-1:DATA_WIDHT*127]}),
            .Valid_Out(Max_Valid_Out)
        );


    Convo_Layer6 #(
        .DATA_WIDHT(DATA_WIDHT),
        .IMG_WIDHT(IMG_WIDHT),
        .IMG_HEIGHT(IMG_HEIGHT)
    )
        convo (
            .Data_In(Data_In),
            .Valid_In(Valid_In),
            .clk(clk),
            .rst(rst),
            .Data_Out(Convo3_Data_Out),
            .Valid_Out(Convo_Valid_Out)
        );

    
    Line_Buffer #(
        .LENGHT(139),
        .DATA_WIDTH(32)
    )
        lb[127:0] (
            .clk(clk),
            .rst(rst),
            .Valid_In(Convo_Valid_Out),
            .Data_In({Convo3_Data_Out[DATA_WIDHT-1:0], Convo3_Data_Out[DATA_WIDHT*2-1:DATA_WIDHT],Convo3_Data_Out[DATA_WIDHT*3-1:DATA_WIDHT*2],Convo3_Data_Out[DATA_WIDHT*4-1:DATA_WIDHT*3],Convo3_Data_Out[DATA_WIDHT*5-1:DATA_WIDHT*4],Convo3_Data_Out[DATA_WIDHT*6-1:DATA_WIDHT*5],Convo3_Data_Out[DATA_WIDHT*7-1:DATA_WIDHT*6],Convo3_Data_Out[DATA_WIDHT*8-1:DATA_WIDHT*7],Convo3_Data_Out[DATA_WIDHT*9-1:DATA_WIDHT*8],Convo3_Data_Out[DATA_WIDHT*10-1:DATA_WIDHT*9],Convo3_Data_Out[DATA_WIDHT*11-1:DATA_WIDHT*10],Convo3_Data_Out[DATA_WIDHT*12-1:DATA_WIDHT*11],Convo3_Data_Out[DATA_WIDHT*13-1:DATA_WIDHT*12],Convo3_Data_Out[DATA_WIDHT*14-1:DATA_WIDHT*13],Convo3_Data_Out[DATA_WIDHT*15-1:DATA_WIDHT*14],Convo3_Data_Out[DATA_WIDHT*16-1:DATA_WIDHT*15],Convo3_Data_Out[DATA_WIDHT*17-1:DATA_WIDHT*16],Convo3_Data_Out[DATA_WIDHT*18-1:DATA_WIDHT*17],Convo3_Data_Out[DATA_WIDHT*19-1:DATA_WIDHT*18],Convo3_Data_Out[DATA_WIDHT*20-1:DATA_WIDHT*19],Convo3_Data_Out[DATA_WIDHT*21-1:DATA_WIDHT*20],Convo3_Data_Out[DATA_WIDHT*22-1:DATA_WIDHT*21],Convo3_Data_Out[DATA_WIDHT*23-1:DATA_WIDHT*22],Convo3_Data_Out[DATA_WIDHT*24-1:DATA_WIDHT*23],Convo3_Data_Out[DATA_WIDHT*25-1:DATA_WIDHT*24],Convo3_Data_Out[DATA_WIDHT*26-1:DATA_WIDHT*25],Convo3_Data_Out[DATA_WIDHT*27-1:DATA_WIDHT*26],Convo3_Data_Out[DATA_WIDHT*28-1:DATA_WIDHT*27],Convo3_Data_Out[DATA_WIDHT*29-1:DATA_WIDHT*28],Convo3_Data_Out[DATA_WIDHT*30-1:DATA_WIDHT*29],Convo3_Data_Out[DATA_WIDHT*31-1:DATA_WIDHT*30],Convo3_Data_Out[DATA_WIDHT*32-1:DATA_WIDHT*31],Convo3_Data_Out[DATA_WIDHT*33-1:DATA_WIDHT*32],Convo3_Data_Out[DATA_WIDHT*34-1:DATA_WIDHT*33],Convo3_Data_Out[DATA_WIDHT*35-1:DATA_WIDHT*34],Convo3_Data_Out[DATA_WIDHT*36-1:DATA_WIDHT*35],Convo3_Data_Out[DATA_WIDHT*37-1:DATA_WIDHT*36],Convo3_Data_Out[DATA_WIDHT*38-1:DATA_WIDHT*37],Convo3_Data_Out[DATA_WIDHT*39-1:DATA_WIDHT*38],Convo3_Data_Out[DATA_WIDHT*40-1:DATA_WIDHT*39],Convo3_Data_Out[DATA_WIDHT*41-1:DATA_WIDHT*40],Convo3_Data_Out[DATA_WIDHT*42-1:DATA_WIDHT*41],Convo3_Data_Out[DATA_WIDHT*43-1:DATA_WIDHT*42],Convo3_Data_Out[DATA_WIDHT*44-1:DATA_WIDHT*43],Convo3_Data_Out[DATA_WIDHT*45-1:DATA_WIDHT*44],Convo3_Data_Out[DATA_WIDHT*46-1:DATA_WIDHT*45],Convo3_Data_Out[DATA_WIDHT*47-1:DATA_WIDHT*46],Convo3_Data_Out[DATA_WIDHT*48-1:DATA_WIDHT*47],Convo3_Data_Out[DATA_WIDHT*49-1:DATA_WIDHT*48],Convo3_Data_Out[DATA_WIDHT*50-1:DATA_WIDHT*49],Convo3_Data_Out[DATA_WIDHT*51-1:DATA_WIDHT*50],Convo3_Data_Out[DATA_WIDHT*52-1:DATA_WIDHT*51],Convo3_Data_Out[DATA_WIDHT*53-1:DATA_WIDHT*52],Convo3_Data_Out[DATA_WIDHT*54-1:DATA_WIDHT*53],Convo3_Data_Out[DATA_WIDHT*55-1:DATA_WIDHT*54],Convo3_Data_Out[DATA_WIDHT*56-1:DATA_WIDHT*55],Convo3_Data_Out[DATA_WIDHT*57-1:DATA_WIDHT*56],Convo3_Data_Out[DATA_WIDHT*58-1:DATA_WIDHT*57],Convo3_Data_Out[DATA_WIDHT*59-1:DATA_WIDHT*58],Convo3_Data_Out[DATA_WIDHT*60-1:DATA_WIDHT*59],Convo3_Data_Out[DATA_WIDHT*61-1:DATA_WIDHT*60],Convo3_Data_Out[DATA_WIDHT*62-1:DATA_WIDHT*61],Convo3_Data_Out[DATA_WIDHT*63-1:DATA_WIDHT*62],Convo3_Data_Out[DATA_WIDHT*64-1:DATA_WIDHT*63],Convo3_Data_Out[DATA_WIDHT*65-1:DATA_WIDHT*64],Convo3_Data_Out[DATA_WIDHT*66-1:DATA_WIDHT*65],Convo3_Data_Out[DATA_WIDHT*67-1:DATA_WIDHT*66],Convo3_Data_Out[DATA_WIDHT*68-1:DATA_WIDHT*67],Convo3_Data_Out[DATA_WIDHT*69-1:DATA_WIDHT*68],Convo3_Data_Out[DATA_WIDHT*70-1:DATA_WIDHT*69],Convo3_Data_Out[DATA_WIDHT*71-1:DATA_WIDHT*70],Convo3_Data_Out[DATA_WIDHT*72-1:DATA_WIDHT*71],Convo3_Data_Out[DATA_WIDHT*73-1:DATA_WIDHT*72],Convo3_Data_Out[DATA_WIDHT*74-1:DATA_WIDHT*73],Convo3_Data_Out[DATA_WIDHT*75-1:DATA_WIDHT*74],Convo3_Data_Out[DATA_WIDHT*76-1:DATA_WIDHT*75],Convo3_Data_Out[DATA_WIDHT*77-1:DATA_WIDHT*76],Convo3_Data_Out[DATA_WIDHT*78-1:DATA_WIDHT*77],Convo3_Data_Out[DATA_WIDHT*79-1:DATA_WIDHT*78],Convo3_Data_Out[DATA_WIDHT*80-1:DATA_WIDHT*79],Convo3_Data_Out[DATA_WIDHT*81-1:DATA_WIDHT*80],Convo3_Data_Out[DATA_WIDHT*82-1:DATA_WIDHT*81],Convo3_Data_Out[DATA_WIDHT*83-1:DATA_WIDHT*82],Convo3_Data_Out[DATA_WIDHT*84-1:DATA_WIDHT*83],Convo3_Data_Out[DATA_WIDHT*85-1:DATA_WIDHT*84],Convo3_Data_Out[DATA_WIDHT*86-1:DATA_WIDHT*85],Convo3_Data_Out[DATA_WIDHT*87-1:DATA_WIDHT*86],Convo3_Data_Out[DATA_WIDHT*88-1:DATA_WIDHT*87],Convo3_Data_Out[DATA_WIDHT*89-1:DATA_WIDHT*88],Convo3_Data_Out[DATA_WIDHT*90-1:DATA_WIDHT*89],Convo3_Data_Out[DATA_WIDHT*91-1:DATA_WIDHT*90],Convo3_Data_Out[DATA_WIDHT*92-1:DATA_WIDHT*91],Convo3_Data_Out[DATA_WIDHT*93-1:DATA_WIDHT*92],Convo3_Data_Out[DATA_WIDHT*94-1:DATA_WIDHT*93],Convo3_Data_Out[DATA_WIDHT*95-1:DATA_WIDHT*94],Convo3_Data_Out[DATA_WIDHT*96-1:DATA_WIDHT*95],Convo3_Data_Out[DATA_WIDHT*97-1:DATA_WIDHT*96],Convo3_Data_Out[DATA_WIDHT*98-1:DATA_WIDHT*97],Convo3_Data_Out[DATA_WIDHT*99-1:DATA_WIDHT*98],Convo3_Data_Out[DATA_WIDHT*100-1:DATA_WIDHT*99],Convo3_Data_Out[DATA_WIDHT*101-1:DATA_WIDHT*100],Convo3_Data_Out[DATA_WIDHT*102-1:DATA_WIDHT*101],Convo3_Data_Out[DATA_WIDHT*103-1:DATA_WIDHT*102],Convo3_Data_Out[DATA_WIDHT*104-1:DATA_WIDHT*103],Convo3_Data_Out[DATA_WIDHT*105-1:DATA_WIDHT*104],Convo3_Data_Out[DATA_WIDHT*106-1:DATA_WIDHT*105],Convo3_Data_Out[DATA_WIDHT*107-1:DATA_WIDHT*106],Convo3_Data_Out[DATA_WIDHT*108-1:DATA_WIDHT*107],Convo3_Data_Out[DATA_WIDHT*109-1:DATA_WIDHT*108],Convo3_Data_Out[DATA_WIDHT*110-1:DATA_WIDHT*109],Convo3_Data_Out[DATA_WIDHT*111-1:DATA_WIDHT*110],Convo3_Data_Out[DATA_WIDHT*112-1:DATA_WIDHT*111],Convo3_Data_Out[DATA_WIDHT*113-1:DATA_WIDHT*112],Convo3_Data_Out[DATA_WIDHT*114-1:DATA_WIDHT*113],Convo3_Data_Out[DATA_WIDHT*115-1:DATA_WIDHT*114],Convo3_Data_Out[DATA_WIDHT*116-1:DATA_WIDHT*115],Convo3_Data_Out[DATA_WIDHT*117-1:DATA_WIDHT*116],Convo3_Data_Out[DATA_WIDHT*118-1:DATA_WIDHT*117],Convo3_Data_Out[DATA_WIDHT*119-1:DATA_WIDHT*118],Convo3_Data_Out[DATA_WIDHT*120-1:DATA_WIDHT*119],Convo3_Data_Out[DATA_WIDHT*121-1:DATA_WIDHT*120],Convo3_Data_Out[DATA_WIDHT*122-1:DATA_WIDHT*121],Convo3_Data_Out[DATA_WIDHT*123-1:DATA_WIDHT*122],Convo3_Data_Out[DATA_WIDHT*124-1:DATA_WIDHT*123],Convo3_Data_Out[DATA_WIDHT*125-1:DATA_WIDHT*124],Convo3_Data_Out[DATA_WIDHT*126-1:DATA_WIDHT*125],Convo3_Data_Out[DATA_WIDHT*127-1:DATA_WIDHT*126],Convo3_Data_Out[DATA_WIDHT*128-1:DATA_WIDHT*127]}),
            .Valid_Out(lb_Valid_Out),
            .Data_Out({lb_Data_Out[DATA_WIDHT-1:0], lb_Data_Out[DATA_WIDHT*2-1:DATA_WIDHT],lb_Data_Out[DATA_WIDHT*3-1:DATA_WIDHT*2],lb_Data_Out[DATA_WIDHT*4-1:DATA_WIDHT*3],lb_Data_Out[DATA_WIDHT*5-1:DATA_WIDHT*4],lb_Data_Out[DATA_WIDHT*6-1:DATA_WIDHT*5],lb_Data_Out[DATA_WIDHT*7-1:DATA_WIDHT*6],lb_Data_Out[DATA_WIDHT*8-1:DATA_WIDHT*7],lb_Data_Out[DATA_WIDHT*9-1:DATA_WIDHT*8],lb_Data_Out[DATA_WIDHT*10-1:DATA_WIDHT*9],lb_Data_Out[DATA_WIDHT*11-1:DATA_WIDHT*10],lb_Data_Out[DATA_WIDHT*12-1:DATA_WIDHT*11],lb_Data_Out[DATA_WIDHT*13-1:DATA_WIDHT*12],lb_Data_Out[DATA_WIDHT*14-1:DATA_WIDHT*13],lb_Data_Out[DATA_WIDHT*15-1:DATA_WIDHT*14],lb_Data_Out[DATA_WIDHT*16-1:DATA_WIDHT*15],lb_Data_Out[DATA_WIDHT*17-1:DATA_WIDHT*16],lb_Data_Out[DATA_WIDHT*18-1:DATA_WIDHT*17],lb_Data_Out[DATA_WIDHT*19-1:DATA_WIDHT*18],lb_Data_Out[DATA_WIDHT*20-1:DATA_WIDHT*19],lb_Data_Out[DATA_WIDHT*21-1:DATA_WIDHT*20],lb_Data_Out[DATA_WIDHT*22-1:DATA_WIDHT*21],lb_Data_Out[DATA_WIDHT*23-1:DATA_WIDHT*22],lb_Data_Out[DATA_WIDHT*24-1:DATA_WIDHT*23],lb_Data_Out[DATA_WIDHT*25-1:DATA_WIDHT*24],lb_Data_Out[DATA_WIDHT*26-1:DATA_WIDHT*25],lb_Data_Out[DATA_WIDHT*27-1:DATA_WIDHT*26],lb_Data_Out[DATA_WIDHT*28-1:DATA_WIDHT*27],lb_Data_Out[DATA_WIDHT*29-1:DATA_WIDHT*28],lb_Data_Out[DATA_WIDHT*30-1:DATA_WIDHT*29],lb_Data_Out[DATA_WIDHT*31-1:DATA_WIDHT*30],lb_Data_Out[DATA_WIDHT*32-1:DATA_WIDHT*31],lb_Data_Out[DATA_WIDHT*33-1:DATA_WIDHT*32],lb_Data_Out[DATA_WIDHT*34-1:DATA_WIDHT*33],lb_Data_Out[DATA_WIDHT*35-1:DATA_WIDHT*34],lb_Data_Out[DATA_WIDHT*36-1:DATA_WIDHT*35],lb_Data_Out[DATA_WIDHT*37-1:DATA_WIDHT*36],lb_Data_Out[DATA_WIDHT*38-1:DATA_WIDHT*37],lb_Data_Out[DATA_WIDHT*39-1:DATA_WIDHT*38],lb_Data_Out[DATA_WIDHT*40-1:DATA_WIDHT*39],lb_Data_Out[DATA_WIDHT*41-1:DATA_WIDHT*40],lb_Data_Out[DATA_WIDHT*42-1:DATA_WIDHT*41],lb_Data_Out[DATA_WIDHT*43-1:DATA_WIDHT*42],lb_Data_Out[DATA_WIDHT*44-1:DATA_WIDHT*43],lb_Data_Out[DATA_WIDHT*45-1:DATA_WIDHT*44],lb_Data_Out[DATA_WIDHT*46-1:DATA_WIDHT*45],lb_Data_Out[DATA_WIDHT*47-1:DATA_WIDHT*46],lb_Data_Out[DATA_WIDHT*48-1:DATA_WIDHT*47],lb_Data_Out[DATA_WIDHT*49-1:DATA_WIDHT*48],lb_Data_Out[DATA_WIDHT*50-1:DATA_WIDHT*49],lb_Data_Out[DATA_WIDHT*51-1:DATA_WIDHT*50],lb_Data_Out[DATA_WIDHT*52-1:DATA_WIDHT*51],lb_Data_Out[DATA_WIDHT*53-1:DATA_WIDHT*52],lb_Data_Out[DATA_WIDHT*54-1:DATA_WIDHT*53],lb_Data_Out[DATA_WIDHT*55-1:DATA_WIDHT*54],lb_Data_Out[DATA_WIDHT*56-1:DATA_WIDHT*55],lb_Data_Out[DATA_WIDHT*57-1:DATA_WIDHT*56],lb_Data_Out[DATA_WIDHT*58-1:DATA_WIDHT*57],lb_Data_Out[DATA_WIDHT*59-1:DATA_WIDHT*58],lb_Data_Out[DATA_WIDHT*60-1:DATA_WIDHT*59],lb_Data_Out[DATA_WIDHT*61-1:DATA_WIDHT*60],lb_Data_Out[DATA_WIDHT*62-1:DATA_WIDHT*61],lb_Data_Out[DATA_WIDHT*63-1:DATA_WIDHT*62],lb_Data_Out[DATA_WIDHT*64-1:DATA_WIDHT*63],lb_Data_Out[DATA_WIDHT*65-1:DATA_WIDHT*64],lb_Data_Out[DATA_WIDHT*66-1:DATA_WIDHT*65],lb_Data_Out[DATA_WIDHT*67-1:DATA_WIDHT*66],lb_Data_Out[DATA_WIDHT*68-1:DATA_WIDHT*67],lb_Data_Out[DATA_WIDHT*69-1:DATA_WIDHT*68],lb_Data_Out[DATA_WIDHT*70-1:DATA_WIDHT*69],lb_Data_Out[DATA_WIDHT*71-1:DATA_WIDHT*70],lb_Data_Out[DATA_WIDHT*72-1:DATA_WIDHT*71],lb_Data_Out[DATA_WIDHT*73-1:DATA_WIDHT*72],lb_Data_Out[DATA_WIDHT*74-1:DATA_WIDHT*73],lb_Data_Out[DATA_WIDHT*75-1:DATA_WIDHT*74],lb_Data_Out[DATA_WIDHT*76-1:DATA_WIDHT*75],lb_Data_Out[DATA_WIDHT*77-1:DATA_WIDHT*76],lb_Data_Out[DATA_WIDHT*78-1:DATA_WIDHT*77],lb_Data_Out[DATA_WIDHT*79-1:DATA_WIDHT*78],lb_Data_Out[DATA_WIDHT*80-1:DATA_WIDHT*79],lb_Data_Out[DATA_WIDHT*81-1:DATA_WIDHT*80],lb_Data_Out[DATA_WIDHT*82-1:DATA_WIDHT*81],lb_Data_Out[DATA_WIDHT*83-1:DATA_WIDHT*82],lb_Data_Out[DATA_WIDHT*84-1:DATA_WIDHT*83],lb_Data_Out[DATA_WIDHT*85-1:DATA_WIDHT*84],lb_Data_Out[DATA_WIDHT*86-1:DATA_WIDHT*85],lb_Data_Out[DATA_WIDHT*87-1:DATA_WIDHT*86],lb_Data_Out[DATA_WIDHT*88-1:DATA_WIDHT*87],lb_Data_Out[DATA_WIDHT*89-1:DATA_WIDHT*88],lb_Data_Out[DATA_WIDHT*90-1:DATA_WIDHT*89],lb_Data_Out[DATA_WIDHT*91-1:DATA_WIDHT*90],lb_Data_Out[DATA_WIDHT*92-1:DATA_WIDHT*91],lb_Data_Out[DATA_WIDHT*93-1:DATA_WIDHT*92],lb_Data_Out[DATA_WIDHT*94-1:DATA_WIDHT*93],lb_Data_Out[DATA_WIDHT*95-1:DATA_WIDHT*94],lb_Data_Out[DATA_WIDHT*96-1:DATA_WIDHT*95],lb_Data_Out[DATA_WIDHT*97-1:DATA_WIDHT*96],lb_Data_Out[DATA_WIDHT*98-1:DATA_WIDHT*97],lb_Data_Out[DATA_WIDHT*99-1:DATA_WIDHT*98],lb_Data_Out[DATA_WIDHT*100-1:DATA_WIDHT*99],lb_Data_Out[DATA_WIDHT*101-1:DATA_WIDHT*100],lb_Data_Out[DATA_WIDHT*102-1:DATA_WIDHT*101],lb_Data_Out[DATA_WIDHT*103-1:DATA_WIDHT*102],lb_Data_Out[DATA_WIDHT*104-1:DATA_WIDHT*103],lb_Data_Out[DATA_WIDHT*105-1:DATA_WIDHT*104],lb_Data_Out[DATA_WIDHT*106-1:DATA_WIDHT*105],lb_Data_Out[DATA_WIDHT*107-1:DATA_WIDHT*106],lb_Data_Out[DATA_WIDHT*108-1:DATA_WIDHT*107],lb_Data_Out[DATA_WIDHT*109-1:DATA_WIDHT*108],lb_Data_Out[DATA_WIDHT*110-1:DATA_WIDHT*109],lb_Data_Out[DATA_WIDHT*111-1:DATA_WIDHT*110],lb_Data_Out[DATA_WIDHT*112-1:DATA_WIDHT*111],lb_Data_Out[DATA_WIDHT*113-1:DATA_WIDHT*112],lb_Data_Out[DATA_WIDHT*114-1:DATA_WIDHT*113],lb_Data_Out[DATA_WIDHT*115-1:DATA_WIDHT*114],lb_Data_Out[DATA_WIDHT*116-1:DATA_WIDHT*115],lb_Data_Out[DATA_WIDHT*117-1:DATA_WIDHT*116],lb_Data_Out[DATA_WIDHT*118-1:DATA_WIDHT*117],lb_Data_Out[DATA_WIDHT*119-1:DATA_WIDHT*118],lb_Data_Out[DATA_WIDHT*120-1:DATA_WIDHT*119],lb_Data_Out[DATA_WIDHT*121-1:DATA_WIDHT*120],lb_Data_Out[DATA_WIDHT*122-1:DATA_WIDHT*121],lb_Data_Out[DATA_WIDHT*123-1:DATA_WIDHT*122],lb_Data_Out[DATA_WIDHT*124-1:DATA_WIDHT*123],lb_Data_Out[DATA_WIDHT*125-1:DATA_WIDHT*124],lb_Data_Out[DATA_WIDHT*126-1:DATA_WIDHT*125],lb_Data_Out[DATA_WIDHT*127-1:DATA_WIDHT*126],lb_Data_Out[DATA_WIDHT*128-1:DATA_WIDHT*127]})
        );


    FP_Adder adder[127:0] (
        .Data_A({Max_Data_Out[DATA_WIDHT-1:0], Max_Data_Out[DATA_WIDHT*2-1:DATA_WIDHT],Max_Data_Out[DATA_WIDHT*3-1:DATA_WIDHT*2],Max_Data_Out[DATA_WIDHT*4-1:DATA_WIDHT*3],Max_Data_Out[DATA_WIDHT*5-1:DATA_WIDHT*4],Max_Data_Out[DATA_WIDHT*6-1:DATA_WIDHT*5],Max_Data_Out[DATA_WIDHT*7-1:DATA_WIDHT*6],Max_Data_Out[DATA_WIDHT*8-1:DATA_WIDHT*7],Max_Data_Out[DATA_WIDHT*9-1:DATA_WIDHT*8],Max_Data_Out[DATA_WIDHT*10-1:DATA_WIDHT*9],Max_Data_Out[DATA_WIDHT*11-1:DATA_WIDHT*10],Max_Data_Out[DATA_WIDHT*12-1:DATA_WIDHT*11],Max_Data_Out[DATA_WIDHT*13-1:DATA_WIDHT*12],Max_Data_Out[DATA_WIDHT*14-1:DATA_WIDHT*13],Max_Data_Out[DATA_WIDHT*15-1:DATA_WIDHT*14],Max_Data_Out[DATA_WIDHT*16-1:DATA_WIDHT*15],Max_Data_Out[DATA_WIDHT*17-1:DATA_WIDHT*16],Max_Data_Out[DATA_WIDHT*18-1:DATA_WIDHT*17],Max_Data_Out[DATA_WIDHT*19-1:DATA_WIDHT*18],Max_Data_Out[DATA_WIDHT*20-1:DATA_WIDHT*19],Max_Data_Out[DATA_WIDHT*21-1:DATA_WIDHT*20],Max_Data_Out[DATA_WIDHT*22-1:DATA_WIDHT*21],Max_Data_Out[DATA_WIDHT*23-1:DATA_WIDHT*22],Max_Data_Out[DATA_WIDHT*24-1:DATA_WIDHT*23],Max_Data_Out[DATA_WIDHT*25-1:DATA_WIDHT*24],Max_Data_Out[DATA_WIDHT*26-1:DATA_WIDHT*25],Max_Data_Out[DATA_WIDHT*27-1:DATA_WIDHT*26],Max_Data_Out[DATA_WIDHT*28-1:DATA_WIDHT*27],Max_Data_Out[DATA_WIDHT*29-1:DATA_WIDHT*28],Max_Data_Out[DATA_WIDHT*30-1:DATA_WIDHT*29],Max_Data_Out[DATA_WIDHT*31-1:DATA_WIDHT*30],Max_Data_Out[DATA_WIDHT*32-1:DATA_WIDHT*31],Max_Data_Out[DATA_WIDHT*33-1:DATA_WIDHT*32],Max_Data_Out[DATA_WIDHT*34-1:DATA_WIDHT*33],Max_Data_Out[DATA_WIDHT*35-1:DATA_WIDHT*34],Max_Data_Out[DATA_WIDHT*36-1:DATA_WIDHT*35],Max_Data_Out[DATA_WIDHT*37-1:DATA_WIDHT*36],Max_Data_Out[DATA_WIDHT*38-1:DATA_WIDHT*37],Max_Data_Out[DATA_WIDHT*39-1:DATA_WIDHT*38],Max_Data_Out[DATA_WIDHT*40-1:DATA_WIDHT*39],Max_Data_Out[DATA_WIDHT*41-1:DATA_WIDHT*40],Max_Data_Out[DATA_WIDHT*42-1:DATA_WIDHT*41],Max_Data_Out[DATA_WIDHT*43-1:DATA_WIDHT*42],Max_Data_Out[DATA_WIDHT*44-1:DATA_WIDHT*43],Max_Data_Out[DATA_WIDHT*45-1:DATA_WIDHT*44],Max_Data_Out[DATA_WIDHT*46-1:DATA_WIDHT*45],Max_Data_Out[DATA_WIDHT*47-1:DATA_WIDHT*46],Max_Data_Out[DATA_WIDHT*48-1:DATA_WIDHT*47],Max_Data_Out[DATA_WIDHT*49-1:DATA_WIDHT*48],Max_Data_Out[DATA_WIDHT*50-1:DATA_WIDHT*49],Max_Data_Out[DATA_WIDHT*51-1:DATA_WIDHT*50],Max_Data_Out[DATA_WIDHT*52-1:DATA_WIDHT*51],Max_Data_Out[DATA_WIDHT*53-1:DATA_WIDHT*52],Max_Data_Out[DATA_WIDHT*54-1:DATA_WIDHT*53],Max_Data_Out[DATA_WIDHT*55-1:DATA_WIDHT*54],Max_Data_Out[DATA_WIDHT*56-1:DATA_WIDHT*55],Max_Data_Out[DATA_WIDHT*57-1:DATA_WIDHT*56],Max_Data_Out[DATA_WIDHT*58-1:DATA_WIDHT*57],Max_Data_Out[DATA_WIDHT*59-1:DATA_WIDHT*58],Max_Data_Out[DATA_WIDHT*60-1:DATA_WIDHT*59],Max_Data_Out[DATA_WIDHT*61-1:DATA_WIDHT*60],Max_Data_Out[DATA_WIDHT*62-1:DATA_WIDHT*61],Max_Data_Out[DATA_WIDHT*63-1:DATA_WIDHT*62],Max_Data_Out[DATA_WIDHT*64-1:DATA_WIDHT*63],Max_Data_Out[DATA_WIDHT*65-1:DATA_WIDHT*64],Max_Data_Out[DATA_WIDHT*66-1:DATA_WIDHT*65],Max_Data_Out[DATA_WIDHT*67-1:DATA_WIDHT*66],Max_Data_Out[DATA_WIDHT*68-1:DATA_WIDHT*67],Max_Data_Out[DATA_WIDHT*69-1:DATA_WIDHT*68],Max_Data_Out[DATA_WIDHT*70-1:DATA_WIDHT*69],Max_Data_Out[DATA_WIDHT*71-1:DATA_WIDHT*70],Max_Data_Out[DATA_WIDHT*72-1:DATA_WIDHT*71],Max_Data_Out[DATA_WIDHT*73-1:DATA_WIDHT*72],Max_Data_Out[DATA_WIDHT*74-1:DATA_WIDHT*73],Max_Data_Out[DATA_WIDHT*75-1:DATA_WIDHT*74],Max_Data_Out[DATA_WIDHT*76-1:DATA_WIDHT*75],Max_Data_Out[DATA_WIDHT*77-1:DATA_WIDHT*76],Max_Data_Out[DATA_WIDHT*78-1:DATA_WIDHT*77],Max_Data_Out[DATA_WIDHT*79-1:DATA_WIDHT*78],Max_Data_Out[DATA_WIDHT*80-1:DATA_WIDHT*79],Max_Data_Out[DATA_WIDHT*81-1:DATA_WIDHT*80],Max_Data_Out[DATA_WIDHT*82-1:DATA_WIDHT*81],Max_Data_Out[DATA_WIDHT*83-1:DATA_WIDHT*82],Max_Data_Out[DATA_WIDHT*84-1:DATA_WIDHT*83],Max_Data_Out[DATA_WIDHT*85-1:DATA_WIDHT*84],Max_Data_Out[DATA_WIDHT*86-1:DATA_WIDHT*85],Max_Data_Out[DATA_WIDHT*87-1:DATA_WIDHT*86],Max_Data_Out[DATA_WIDHT*88-1:DATA_WIDHT*87],Max_Data_Out[DATA_WIDHT*89-1:DATA_WIDHT*88],Max_Data_Out[DATA_WIDHT*90-1:DATA_WIDHT*89],Max_Data_Out[DATA_WIDHT*91-1:DATA_WIDHT*90],Max_Data_Out[DATA_WIDHT*92-1:DATA_WIDHT*91],Max_Data_Out[DATA_WIDHT*93-1:DATA_WIDHT*92],Max_Data_Out[DATA_WIDHT*94-1:DATA_WIDHT*93],Max_Data_Out[DATA_WIDHT*95-1:DATA_WIDHT*94],Max_Data_Out[DATA_WIDHT*96-1:DATA_WIDHT*95],Max_Data_Out[DATA_WIDHT*97-1:DATA_WIDHT*96],Max_Data_Out[DATA_WIDHT*98-1:DATA_WIDHT*97],Max_Data_Out[DATA_WIDHT*99-1:DATA_WIDHT*98],Max_Data_Out[DATA_WIDHT*100-1:DATA_WIDHT*99],Max_Data_Out[DATA_WIDHT*101-1:DATA_WIDHT*100],Max_Data_Out[DATA_WIDHT*102-1:DATA_WIDHT*101],Max_Data_Out[DATA_WIDHT*103-1:DATA_WIDHT*102],Max_Data_Out[DATA_WIDHT*104-1:DATA_WIDHT*103],Max_Data_Out[DATA_WIDHT*105-1:DATA_WIDHT*104],Max_Data_Out[DATA_WIDHT*106-1:DATA_WIDHT*105],Max_Data_Out[DATA_WIDHT*107-1:DATA_WIDHT*106],Max_Data_Out[DATA_WIDHT*108-1:DATA_WIDHT*107],Max_Data_Out[DATA_WIDHT*109-1:DATA_WIDHT*108],Max_Data_Out[DATA_WIDHT*110-1:DATA_WIDHT*109],Max_Data_Out[DATA_WIDHT*111-1:DATA_WIDHT*110],Max_Data_Out[DATA_WIDHT*112-1:DATA_WIDHT*111],Max_Data_Out[DATA_WIDHT*113-1:DATA_WIDHT*112],Max_Data_Out[DATA_WIDHT*114-1:DATA_WIDHT*113],Max_Data_Out[DATA_WIDHT*115-1:DATA_WIDHT*114],Max_Data_Out[DATA_WIDHT*116-1:DATA_WIDHT*115],Max_Data_Out[DATA_WIDHT*117-1:DATA_WIDHT*116],Max_Data_Out[DATA_WIDHT*118-1:DATA_WIDHT*117],Max_Data_Out[DATA_WIDHT*119-1:DATA_WIDHT*118],Max_Data_Out[DATA_WIDHT*120-1:DATA_WIDHT*119],Max_Data_Out[DATA_WIDHT*121-1:DATA_WIDHT*120],Max_Data_Out[DATA_WIDHT*122-1:DATA_WIDHT*121],Max_Data_Out[DATA_WIDHT*123-1:DATA_WIDHT*122],Max_Data_Out[DATA_WIDHT*124-1:DATA_WIDHT*123],Max_Data_Out[DATA_WIDHT*125-1:DATA_WIDHT*124],Max_Data_Out[DATA_WIDHT*126-1:DATA_WIDHT*125],Max_Data_Out[DATA_WIDHT*127-1:DATA_WIDHT*126],Max_Data_Out[DATA_WIDHT*128-1:DATA_WIDHT*127]}),
        .Data_B({lb_Data_Out[DATA_WIDHT-1:0], lb_Data_Out[DATA_WIDHT*2-1:DATA_WIDHT],lb_Data_Out[DATA_WIDHT*3-1:DATA_WIDHT*2],lb_Data_Out[DATA_WIDHT*4-1:DATA_WIDHT*3],lb_Data_Out[DATA_WIDHT*5-1:DATA_WIDHT*4],lb_Data_Out[DATA_WIDHT*6-1:DATA_WIDHT*5],lb_Data_Out[DATA_WIDHT*7-1:DATA_WIDHT*6],lb_Data_Out[DATA_WIDHT*8-1:DATA_WIDHT*7],lb_Data_Out[DATA_WIDHT*9-1:DATA_WIDHT*8],lb_Data_Out[DATA_WIDHT*10-1:DATA_WIDHT*9],lb_Data_Out[DATA_WIDHT*11-1:DATA_WIDHT*10],lb_Data_Out[DATA_WIDHT*12-1:DATA_WIDHT*11],lb_Data_Out[DATA_WIDHT*13-1:DATA_WIDHT*12],lb_Data_Out[DATA_WIDHT*14-1:DATA_WIDHT*13],lb_Data_Out[DATA_WIDHT*15-1:DATA_WIDHT*14],lb_Data_Out[DATA_WIDHT*16-1:DATA_WIDHT*15],lb_Data_Out[DATA_WIDHT*17-1:DATA_WIDHT*16],lb_Data_Out[DATA_WIDHT*18-1:DATA_WIDHT*17],lb_Data_Out[DATA_WIDHT*19-1:DATA_WIDHT*18],lb_Data_Out[DATA_WIDHT*20-1:DATA_WIDHT*19],lb_Data_Out[DATA_WIDHT*21-1:DATA_WIDHT*20],lb_Data_Out[DATA_WIDHT*22-1:DATA_WIDHT*21],lb_Data_Out[DATA_WIDHT*23-1:DATA_WIDHT*22],lb_Data_Out[DATA_WIDHT*24-1:DATA_WIDHT*23],lb_Data_Out[DATA_WIDHT*25-1:DATA_WIDHT*24],lb_Data_Out[DATA_WIDHT*26-1:DATA_WIDHT*25],lb_Data_Out[DATA_WIDHT*27-1:DATA_WIDHT*26],lb_Data_Out[DATA_WIDHT*28-1:DATA_WIDHT*27],lb_Data_Out[DATA_WIDHT*29-1:DATA_WIDHT*28],lb_Data_Out[DATA_WIDHT*30-1:DATA_WIDHT*29],lb_Data_Out[DATA_WIDHT*31-1:DATA_WIDHT*30],lb_Data_Out[DATA_WIDHT*32-1:DATA_WIDHT*31],lb_Data_Out[DATA_WIDHT*33-1:DATA_WIDHT*32],lb_Data_Out[DATA_WIDHT*34-1:DATA_WIDHT*33],lb_Data_Out[DATA_WIDHT*35-1:DATA_WIDHT*34],lb_Data_Out[DATA_WIDHT*36-1:DATA_WIDHT*35],lb_Data_Out[DATA_WIDHT*37-1:DATA_WIDHT*36],lb_Data_Out[DATA_WIDHT*38-1:DATA_WIDHT*37],lb_Data_Out[DATA_WIDHT*39-1:DATA_WIDHT*38],lb_Data_Out[DATA_WIDHT*40-1:DATA_WIDHT*39],lb_Data_Out[DATA_WIDHT*41-1:DATA_WIDHT*40],lb_Data_Out[DATA_WIDHT*42-1:DATA_WIDHT*41],lb_Data_Out[DATA_WIDHT*43-1:DATA_WIDHT*42],lb_Data_Out[DATA_WIDHT*44-1:DATA_WIDHT*43],lb_Data_Out[DATA_WIDHT*45-1:DATA_WIDHT*44],lb_Data_Out[DATA_WIDHT*46-1:DATA_WIDHT*45],lb_Data_Out[DATA_WIDHT*47-1:DATA_WIDHT*46],lb_Data_Out[DATA_WIDHT*48-1:DATA_WIDHT*47],lb_Data_Out[DATA_WIDHT*49-1:DATA_WIDHT*48],lb_Data_Out[DATA_WIDHT*50-1:DATA_WIDHT*49],lb_Data_Out[DATA_WIDHT*51-1:DATA_WIDHT*50],lb_Data_Out[DATA_WIDHT*52-1:DATA_WIDHT*51],lb_Data_Out[DATA_WIDHT*53-1:DATA_WIDHT*52],lb_Data_Out[DATA_WIDHT*54-1:DATA_WIDHT*53],lb_Data_Out[DATA_WIDHT*55-1:DATA_WIDHT*54],lb_Data_Out[DATA_WIDHT*56-1:DATA_WIDHT*55],lb_Data_Out[DATA_WIDHT*57-1:DATA_WIDHT*56],lb_Data_Out[DATA_WIDHT*58-1:DATA_WIDHT*57],lb_Data_Out[DATA_WIDHT*59-1:DATA_WIDHT*58],lb_Data_Out[DATA_WIDHT*60-1:DATA_WIDHT*59],lb_Data_Out[DATA_WIDHT*61-1:DATA_WIDHT*60],lb_Data_Out[DATA_WIDHT*62-1:DATA_WIDHT*61],lb_Data_Out[DATA_WIDHT*63-1:DATA_WIDHT*62],lb_Data_Out[DATA_WIDHT*64-1:DATA_WIDHT*63],lb_Data_Out[DATA_WIDHT*65-1:DATA_WIDHT*64],lb_Data_Out[DATA_WIDHT*66-1:DATA_WIDHT*65],lb_Data_Out[DATA_WIDHT*67-1:DATA_WIDHT*66],lb_Data_Out[DATA_WIDHT*68-1:DATA_WIDHT*67],lb_Data_Out[DATA_WIDHT*69-1:DATA_WIDHT*68],lb_Data_Out[DATA_WIDHT*70-1:DATA_WIDHT*69],lb_Data_Out[DATA_WIDHT*71-1:DATA_WIDHT*70],lb_Data_Out[DATA_WIDHT*72-1:DATA_WIDHT*71],lb_Data_Out[DATA_WIDHT*73-1:DATA_WIDHT*72],lb_Data_Out[DATA_WIDHT*74-1:DATA_WIDHT*73],lb_Data_Out[DATA_WIDHT*75-1:DATA_WIDHT*74],lb_Data_Out[DATA_WIDHT*76-1:DATA_WIDHT*75],lb_Data_Out[DATA_WIDHT*77-1:DATA_WIDHT*76],lb_Data_Out[DATA_WIDHT*78-1:DATA_WIDHT*77],lb_Data_Out[DATA_WIDHT*79-1:DATA_WIDHT*78],lb_Data_Out[DATA_WIDHT*80-1:DATA_WIDHT*79],lb_Data_Out[DATA_WIDHT*81-1:DATA_WIDHT*80],lb_Data_Out[DATA_WIDHT*82-1:DATA_WIDHT*81],lb_Data_Out[DATA_WIDHT*83-1:DATA_WIDHT*82],lb_Data_Out[DATA_WIDHT*84-1:DATA_WIDHT*83],lb_Data_Out[DATA_WIDHT*85-1:DATA_WIDHT*84],lb_Data_Out[DATA_WIDHT*86-1:DATA_WIDHT*85],lb_Data_Out[DATA_WIDHT*87-1:DATA_WIDHT*86],lb_Data_Out[DATA_WIDHT*88-1:DATA_WIDHT*87],lb_Data_Out[DATA_WIDHT*89-1:DATA_WIDHT*88],lb_Data_Out[DATA_WIDHT*90-1:DATA_WIDHT*89],lb_Data_Out[DATA_WIDHT*91-1:DATA_WIDHT*90],lb_Data_Out[DATA_WIDHT*92-1:DATA_WIDHT*91],lb_Data_Out[DATA_WIDHT*93-1:DATA_WIDHT*92],lb_Data_Out[DATA_WIDHT*94-1:DATA_WIDHT*93],lb_Data_Out[DATA_WIDHT*95-1:DATA_WIDHT*94],lb_Data_Out[DATA_WIDHT*96-1:DATA_WIDHT*95],lb_Data_Out[DATA_WIDHT*97-1:DATA_WIDHT*96],lb_Data_Out[DATA_WIDHT*98-1:DATA_WIDHT*97],lb_Data_Out[DATA_WIDHT*99-1:DATA_WIDHT*98],lb_Data_Out[DATA_WIDHT*100-1:DATA_WIDHT*99],lb_Data_Out[DATA_WIDHT*101-1:DATA_WIDHT*100],lb_Data_Out[DATA_WIDHT*102-1:DATA_WIDHT*101],lb_Data_Out[DATA_WIDHT*103-1:DATA_WIDHT*102],lb_Data_Out[DATA_WIDHT*104-1:DATA_WIDHT*103],lb_Data_Out[DATA_WIDHT*105-1:DATA_WIDHT*104],lb_Data_Out[DATA_WIDHT*106-1:DATA_WIDHT*105],lb_Data_Out[DATA_WIDHT*107-1:DATA_WIDHT*106],lb_Data_Out[DATA_WIDHT*108-1:DATA_WIDHT*107],lb_Data_Out[DATA_WIDHT*109-1:DATA_WIDHT*108],lb_Data_Out[DATA_WIDHT*110-1:DATA_WIDHT*109],lb_Data_Out[DATA_WIDHT*111-1:DATA_WIDHT*110],lb_Data_Out[DATA_WIDHT*112-1:DATA_WIDHT*111],lb_Data_Out[DATA_WIDHT*113-1:DATA_WIDHT*112],lb_Data_Out[DATA_WIDHT*114-1:DATA_WIDHT*113],lb_Data_Out[DATA_WIDHT*115-1:DATA_WIDHT*114],lb_Data_Out[DATA_WIDHT*116-1:DATA_WIDHT*115],lb_Data_Out[DATA_WIDHT*117-1:DATA_WIDHT*116],lb_Data_Out[DATA_WIDHT*118-1:DATA_WIDHT*117],lb_Data_Out[DATA_WIDHT*119-1:DATA_WIDHT*118],lb_Data_Out[DATA_WIDHT*120-1:DATA_WIDHT*119],lb_Data_Out[DATA_WIDHT*121-1:DATA_WIDHT*120],lb_Data_Out[DATA_WIDHT*122-1:DATA_WIDHT*121],lb_Data_Out[DATA_WIDHT*123-1:DATA_WIDHT*122],lb_Data_Out[DATA_WIDHT*124-1:DATA_WIDHT*123],lb_Data_Out[DATA_WIDHT*125-1:DATA_WIDHT*124],lb_Data_Out[DATA_WIDHT*126-1:DATA_WIDHT*125],lb_Data_Out[DATA_WIDHT*127-1:DATA_WIDHT*126],lb_Data_Out[DATA_WIDHT*128-1:DATA_WIDHT*127]}),
        .Valid_In(add_Valid_In),
        .Mode(1'b0),
        .RMode(2'b0),
        .Data_Out({Data_Out[DATA_WIDHT-1:0], Data_Out[DATA_WIDHT*2-1:DATA_WIDHT],Data_Out[DATA_WIDHT*3-1:DATA_WIDHT*2],Data_Out[DATA_WIDHT*4-1:DATA_WIDHT*3],Data_Out[DATA_WIDHT*5-1:DATA_WIDHT*4],Data_Out[DATA_WIDHT*6-1:DATA_WIDHT*5],Data_Out[DATA_WIDHT*7-1:DATA_WIDHT*6],Data_Out[DATA_WIDHT*8-1:DATA_WIDHT*7],Data_Out[DATA_WIDHT*9-1:DATA_WIDHT*8],Data_Out[DATA_WIDHT*10-1:DATA_WIDHT*9],Data_Out[DATA_WIDHT*11-1:DATA_WIDHT*10],Data_Out[DATA_WIDHT*12-1:DATA_WIDHT*11],Data_Out[DATA_WIDHT*13-1:DATA_WIDHT*12],Data_Out[DATA_WIDHT*14-1:DATA_WIDHT*13],Data_Out[DATA_WIDHT*15-1:DATA_WIDHT*14],Data_Out[DATA_WIDHT*16-1:DATA_WIDHT*15],Data_Out[DATA_WIDHT*17-1:DATA_WIDHT*16],Data_Out[DATA_WIDHT*18-1:DATA_WIDHT*17],Data_Out[DATA_WIDHT*19-1:DATA_WIDHT*18],Data_Out[DATA_WIDHT*20-1:DATA_WIDHT*19],Data_Out[DATA_WIDHT*21-1:DATA_WIDHT*20],Data_Out[DATA_WIDHT*22-1:DATA_WIDHT*21],Data_Out[DATA_WIDHT*23-1:DATA_WIDHT*22],Data_Out[DATA_WIDHT*24-1:DATA_WIDHT*23],Data_Out[DATA_WIDHT*25-1:DATA_WIDHT*24],Data_Out[DATA_WIDHT*26-1:DATA_WIDHT*25],Data_Out[DATA_WIDHT*27-1:DATA_WIDHT*26],Data_Out[DATA_WIDHT*28-1:DATA_WIDHT*27],Data_Out[DATA_WIDHT*29-1:DATA_WIDHT*28],Data_Out[DATA_WIDHT*30-1:DATA_WIDHT*29],Data_Out[DATA_WIDHT*31-1:DATA_WIDHT*30],Data_Out[DATA_WIDHT*32-1:DATA_WIDHT*31],Data_Out[DATA_WIDHT*33-1:DATA_WIDHT*32],Data_Out[DATA_WIDHT*34-1:DATA_WIDHT*33],Data_Out[DATA_WIDHT*35-1:DATA_WIDHT*34],Data_Out[DATA_WIDHT*36-1:DATA_WIDHT*35],Data_Out[DATA_WIDHT*37-1:DATA_WIDHT*36],Data_Out[DATA_WIDHT*38-1:DATA_WIDHT*37],Data_Out[DATA_WIDHT*39-1:DATA_WIDHT*38],Data_Out[DATA_WIDHT*40-1:DATA_WIDHT*39],Data_Out[DATA_WIDHT*41-1:DATA_WIDHT*40],Data_Out[DATA_WIDHT*42-1:DATA_WIDHT*41],Data_Out[DATA_WIDHT*43-1:DATA_WIDHT*42],Data_Out[DATA_WIDHT*44-1:DATA_WIDHT*43],Data_Out[DATA_WIDHT*45-1:DATA_WIDHT*44],Data_Out[DATA_WIDHT*46-1:DATA_WIDHT*45],Data_Out[DATA_WIDHT*47-1:DATA_WIDHT*46],Data_Out[DATA_WIDHT*48-1:DATA_WIDHT*47],Data_Out[DATA_WIDHT*49-1:DATA_WIDHT*48],Data_Out[DATA_WIDHT*50-1:DATA_WIDHT*49],Data_Out[DATA_WIDHT*51-1:DATA_WIDHT*50],Data_Out[DATA_WIDHT*52-1:DATA_WIDHT*51],Data_Out[DATA_WIDHT*53-1:DATA_WIDHT*52],Data_Out[DATA_WIDHT*54-1:DATA_WIDHT*53],Data_Out[DATA_WIDHT*55-1:DATA_WIDHT*54],Data_Out[DATA_WIDHT*56-1:DATA_WIDHT*55],Data_Out[DATA_WIDHT*57-1:DATA_WIDHT*56],Data_Out[DATA_WIDHT*58-1:DATA_WIDHT*57],Data_Out[DATA_WIDHT*59-1:DATA_WIDHT*58],Data_Out[DATA_WIDHT*60-1:DATA_WIDHT*59],Data_Out[DATA_WIDHT*61-1:DATA_WIDHT*60],Data_Out[DATA_WIDHT*62-1:DATA_WIDHT*61],Data_Out[DATA_WIDHT*63-1:DATA_WIDHT*62],Data_Out[DATA_WIDHT*64-1:DATA_WIDHT*63],Data_Out[DATA_WIDHT*65-1:DATA_WIDHT*64],Data_Out[DATA_WIDHT*66-1:DATA_WIDHT*65],Data_Out[DATA_WIDHT*67-1:DATA_WIDHT*66],Data_Out[DATA_WIDHT*68-1:DATA_WIDHT*67],Data_Out[DATA_WIDHT*69-1:DATA_WIDHT*68],Data_Out[DATA_WIDHT*70-1:DATA_WIDHT*69],Data_Out[DATA_WIDHT*71-1:DATA_WIDHT*70],Data_Out[DATA_WIDHT*72-1:DATA_WIDHT*71],Data_Out[DATA_WIDHT*73-1:DATA_WIDHT*72],Data_Out[DATA_WIDHT*74-1:DATA_WIDHT*73],Data_Out[DATA_WIDHT*75-1:DATA_WIDHT*74],Data_Out[DATA_WIDHT*76-1:DATA_WIDHT*75],Data_Out[DATA_WIDHT*77-1:DATA_WIDHT*76],Data_Out[DATA_WIDHT*78-1:DATA_WIDHT*77],Data_Out[DATA_WIDHT*79-1:DATA_WIDHT*78],Data_Out[DATA_WIDHT*80-1:DATA_WIDHT*79],Data_Out[DATA_WIDHT*81-1:DATA_WIDHT*80],Data_Out[DATA_WIDHT*82-1:DATA_WIDHT*81],Data_Out[DATA_WIDHT*83-1:DATA_WIDHT*82],Data_Out[DATA_WIDHT*84-1:DATA_WIDHT*83],Data_Out[DATA_WIDHT*85-1:DATA_WIDHT*84],Data_Out[DATA_WIDHT*86-1:DATA_WIDHT*85],Data_Out[DATA_WIDHT*87-1:DATA_WIDHT*86],Data_Out[DATA_WIDHT*88-1:DATA_WIDHT*87],Data_Out[DATA_WIDHT*89-1:DATA_WIDHT*88],Data_Out[DATA_WIDHT*90-1:DATA_WIDHT*89],Data_Out[DATA_WIDHT*91-1:DATA_WIDHT*90],Data_Out[DATA_WIDHT*92-1:DATA_WIDHT*91],Data_Out[DATA_WIDHT*93-1:DATA_WIDHT*92],Data_Out[DATA_WIDHT*94-1:DATA_WIDHT*93],Data_Out[DATA_WIDHT*95-1:DATA_WIDHT*94],Data_Out[DATA_WIDHT*96-1:DATA_WIDHT*95],Data_Out[DATA_WIDHT*97-1:DATA_WIDHT*96],Data_Out[DATA_WIDHT*98-1:DATA_WIDHT*97],Data_Out[DATA_WIDHT*99-1:DATA_WIDHT*98],Data_Out[DATA_WIDHT*100-1:DATA_WIDHT*99],Data_Out[DATA_WIDHT*101-1:DATA_WIDHT*100],Data_Out[DATA_WIDHT*102-1:DATA_WIDHT*101],Data_Out[DATA_WIDHT*103-1:DATA_WIDHT*102],Data_Out[DATA_WIDHT*104-1:DATA_WIDHT*103],Data_Out[DATA_WIDHT*105-1:DATA_WIDHT*104],Data_Out[DATA_WIDHT*106-1:DATA_WIDHT*105],Data_Out[DATA_WIDHT*107-1:DATA_WIDHT*106],Data_Out[DATA_WIDHT*108-1:DATA_WIDHT*107],Data_Out[DATA_WIDHT*109-1:DATA_WIDHT*108],Data_Out[DATA_WIDHT*110-1:DATA_WIDHT*109],Data_Out[DATA_WIDHT*111-1:DATA_WIDHT*110],Data_Out[DATA_WIDHT*112-1:DATA_WIDHT*111],Data_Out[DATA_WIDHT*113-1:DATA_WIDHT*112],Data_Out[DATA_WIDHT*114-1:DATA_WIDHT*113],Data_Out[DATA_WIDHT*115-1:DATA_WIDHT*114],Data_Out[DATA_WIDHT*116-1:DATA_WIDHT*115],Data_Out[DATA_WIDHT*117-1:DATA_WIDHT*116],Data_Out[DATA_WIDHT*118-1:DATA_WIDHT*117],Data_Out[DATA_WIDHT*119-1:DATA_WIDHT*118],Data_Out[DATA_WIDHT*120-1:DATA_WIDHT*119],Data_Out[DATA_WIDHT*121-1:DATA_WIDHT*120],Data_Out[DATA_WIDHT*122-1:DATA_WIDHT*121],Data_Out[DATA_WIDHT*123-1:DATA_WIDHT*122],Data_Out[DATA_WIDHT*124-1:DATA_WIDHT*123],Data_Out[DATA_WIDHT*125-1:DATA_WIDHT*124],Data_Out[DATA_WIDHT*126-1:DATA_WIDHT*125],Data_Out[DATA_WIDHT*127-1:DATA_WIDHT*126],Data_Out[DATA_WIDHT*128-1:DATA_WIDHT*127]}),
        .Valid_Out(Valid_Out)
    );
    
endmodule