module Depthwise_Part2_Separable_64CHANNEL_Layer5 #(
    parameter DATA_WIDHT = 32, 
    parameter IMG_WIDHT = 44,
    parameter IMG_HEIGHT =44
)
(
    input [DATA_WIDHT*32-1:0] Data_In,
    input clk,
    input rst,
    input Valid_In,
    output [DATA_WIDHT*64-1:0] Data_Out,
    output Valid_Out
);
 	wire [DATA_WIDHT*32-1:0] Data_Out_Kernel1, Data_Out_Kernel2, Data_Out_Kernel3, Data_Out_Kernel4, Data_Out_Kernel5, Data_Out_Kernel6, Data_Out_Kernel7, Data_Out_Kernel8, Data_Out_Kernel9, Data_Out_Kernel10, Data_Out_Kernel11, Data_Out_Kernel12, Data_Out_Kernel13, Data_Out_Kernel14, Data_Out_Kernel15, Data_Out_Kernel16, Data_Out_Kernel17, Data_Out_Kernel18, Data_Out_Kernel19, Data_Out_Kernel20, Data_Out_Kernel21, Data_Out_Kernel22, Data_Out_Kernel23, Data_Out_Kernel24, Data_Out_Kernel25, Data_Out_Kernel26, Data_Out_Kernel27, Data_Out_Kernel28, Data_Out_Kernel29, Data_Out_Kernel30, Data_Out_Kernel31, Data_Out_Kernel32, Data_Out_Kernel33, Data_Out_Kernel34, Data_Out_Kernel35, Data_Out_Kernel36, Data_Out_Kernel37, Data_Out_Kernel38, Data_Out_Kernel39, Data_Out_Kernel40, Data_Out_Kernel41, Data_Out_Kernel42, Data_Out_Kernel43, Data_Out_Kernel44, Data_Out_Kernel45, Data_Out_Kernel46, Data_Out_Kernel47, Data_Out_Kernel48, Data_Out_Kernel49, Data_Out_Kernel50, Data_Out_Kernel51, Data_Out_Kernel52, Data_Out_Kernel53, Data_Out_Kernel54, Data_Out_Kernel55, Data_Out_Kernel56, Data_Out_Kernel57, Data_Out_Kernel58, Data_Out_Kernel59, Data_Out_Kernel60, Data_Out_Kernel61, Data_Out_Kernel62, Data_Out_Kernel63, Data_Out_Kernel64;

	wire[31:0] add_k1_Data_Out, add_k2_Data_Out, add_k3_Data_Out, add_k4_Data_Out, add_k5_Data_Out, add_k6_Data_Out, add_k7_Data_Out, add_k8_Data_Out, add_k9_Data_Out, add_k10_Data_Out, add_k11_Data_Out, add_k12_Data_Out, add_k13_Data_Out, add_k14_Data_Out, add_k15_Data_Out, add_k16_Data_Out, add_k17_Data_Out, add_k18_Data_Out, add_k19_Data_Out, add_k20_Data_Out, add_k21_Data_Out, add_k22_Data_Out, add_k23_Data_Out, add_k24_Data_Out, add_k25_Data_Out, add_k26_Data_Out, add_k27_Data_Out, add_k28_Data_Out, add_k29_Data_Out, add_k30_Data_Out, add_k31_Data_Out, add_k32_Data_Out, add_k33_Data_Out, add_k34_Data_Out, add_k35_Data_Out, add_k36_Data_Out, add_k37_Data_Out, add_k38_Data_Out, add_k39_Data_Out, add_k40_Data_Out, add_k41_Data_Out, add_k42_Data_Out, add_k43_Data_Out, add_k44_Data_Out, add_k45_Data_Out, add_k46_Data_Out, add_k47_Data_Out, add_k48_Data_Out, add_k49_Data_Out, add_k50_Data_Out, add_k51_Data_Out, add_k52_Data_Out, add_k53_Data_Out, add_k54_Data_Out, add_k55_Data_Out, add_k56_Data_Out, add_k57_Data_Out, add_k58_Data_Out, add_k59_Data_Out, add_k60_Data_Out, add_k61_Data_Out, add_k62_Data_Out, add_k63_Data_Out, add_k64_Data_Out;



	wire add_kernel1_Valid_Out, add_kernel2_Valid_Out, add_kernel3_Valid_Out, add_kernel4_Valid_Out, add_kernel5_Valid_Out, add_kernel6_Valid_Out, add_kernel7_Valid_Out, add_kernel8_Valid_Out, add_kernel9_Valid_Out, add_kernel10_Valid_Out, add_kernel11_Valid_Out, add_kernel12_Valid_Out, add_kernel13_Valid_Out, add_kernel14_Valid_Out, add_kernel15_Valid_Out, add_kernel16_Valid_Out, add_kernel17_Valid_Out, add_kernel18_Valid_Out, add_kernel19_Valid_Out, add_kernel20_Valid_Out, add_kernel21_Valid_Out, add_kernel22_Valid_Out, add_kernel23_Valid_Out, add_kernel24_Valid_Out, add_kernel25_Valid_Out, add_kernel26_Valid_Out, add_kernel27_Valid_Out, add_kernel28_Valid_Out, add_kernel29_Valid_Out, add_kernel30_Valid_Out, add_kernel31_Valid_Out, add_kernel32_Valid_Out, add_kernel33_Valid_Out, add_kernel34_Valid_Out, add_kernel35_Valid_Out, add_kernel36_Valid_Out, add_kernel37_Valid_Out, add_kernel38_Valid_Out, add_kernel39_Valid_Out, add_kernel40_Valid_Out, add_kernel41_Valid_Out, add_kernel42_Valid_Out, add_kernel43_Valid_Out, add_kernel44_Valid_Out, add_kernel45_Valid_Out, add_kernel46_Valid_Out, add_kernel47_Valid_Out, add_kernel48_Valid_Out, add_kernel49_Valid_Out, add_kernel50_Valid_Out, add_kernel51_Valid_Out, add_kernel52_Valid_Out, add_kernel53_Valid_Out, add_kernel54_Valid_Out, add_kernel55_Valid_Out, add_kernel56_Valid_Out, add_kernel57_Valid_Out, add_kernel58_Valid_Out, add_kernel59_Valid_Out, add_kernel60_Valid_Out, add_kernel61_Valid_Out, add_kernel62_Valid_Out, add_kernel63_Valid_Out, add_kernel64_Valid_Out;

	wire channel1_Kernel1_Valid_Out, channel2_Kernel1_Valid_Out, channel3_Kernel1_Valid_Out, channel4_Kernel1_Valid_Out, channel5_Kernel1_Valid_Out, channel6_Kernel1_Valid_Out, channel7_Kernel1_Valid_Out, channel8_Kernel1_Valid_Out, channel9_Kernel1_Valid_Out, channel10_Kernel1_Valid_Out, channel11_Kernel1_Valid_Out, channel12_Kernel1_Valid_Out, channel13_Kernel1_Valid_Out, channel14_Kernel1_Valid_Out, channel15_Kernel1_Valid_Out, channel16_Kernel1_Valid_Out, channel17_Kernel1_Valid_Out, channel18_Kernel1_Valid_Out, channel19_Kernel1_Valid_Out, channel20_Kernel1_Valid_Out, channel21_Kernel1_Valid_Out, channel22_Kernel1_Valid_Out, channel23_Kernel1_Valid_Out, channel24_Kernel1_Valid_Out, channel25_Kernel1_Valid_Out, channel26_Kernel1_Valid_Out, channel27_Kernel1_Valid_Out, channel28_Kernel1_Valid_Out, channel29_Kernel1_Valid_Out, channel30_Kernel1_Valid_Out, channel31_Kernel1_Valid_Out, channel32_Kernel1_Valid_Out;

	assign add_kernel1=channel1_Kernel1_Valid_Out & channel2_Kernel1_Valid_Out & channel3_Kernel1_Valid_Out & channel4_Kernel1_Valid_Out & channel5_Kernel1_Valid_Out & channel6_Kernel1_Valid_Out & channel7_Kernel1_Valid_Out & channel8_Kernel1_Valid_Out & channel9_Kernel1_Valid_Out & channel10_Kernel1_Valid_Out & channel11_Kernel1_Valid_Out & channel12_Kernel1_Valid_Out & channel13_Kernel1_Valid_Out & channel14_Kernel1_Valid_Out & channel15_Kernel1_Valid_Out & channel16_Kernel1_Valid_Out & channel17_Kernel1_Valid_Out & channel18_Kernel1_Valid_Out & channel19_Kernel1_Valid_Out & channel20_Kernel1_Valid_Out & channel21_Kernel1_Valid_Out & channel22_Kernel1_Valid_Out & channel23_Kernel1_Valid_Out & channel24_Kernel1_Valid_Out & channel25_Kernel1_Valid_Out & channel26_Kernel1_Valid_Out & channel27_Kernel1_Valid_Out & channel28_Kernel1_Valid_Out & channel29_Kernel1_Valid_Out & channel30_Kernel1_Valid_Out & channel31_Kernel1_Valid_Out & channel32_Kernel1_Valid_Out;

	wire channel1_Kernel2_Valid_Out, channel2_Kernel2_Valid_Out, channel3_Kernel2_Valid_Out, channel4_Kernel2_Valid_Out, channel5_Kernel2_Valid_Out, channel6_Kernel2_Valid_Out, channel7_Kernel2_Valid_Out, channel8_Kernel2_Valid_Out, channel9_Kernel2_Valid_Out, channel10_Kernel2_Valid_Out, channel11_Kernel2_Valid_Out, channel12_Kernel2_Valid_Out, channel13_Kernel2_Valid_Out, channel14_Kernel2_Valid_Out, channel15_Kernel2_Valid_Out, channel16_Kernel2_Valid_Out, channel17_Kernel2_Valid_Out, channel18_Kernel2_Valid_Out, channel19_Kernel2_Valid_Out, channel20_Kernel2_Valid_Out, channel21_Kernel2_Valid_Out, channel22_Kernel2_Valid_Out, channel23_Kernel2_Valid_Out, channel24_Kernel2_Valid_Out, channel25_Kernel2_Valid_Out, channel26_Kernel2_Valid_Out, channel27_Kernel2_Valid_Out, channel28_Kernel2_Valid_Out, channel29_Kernel2_Valid_Out, channel30_Kernel2_Valid_Out, channel31_Kernel2_Valid_Out, channel32_Kernel2_Valid_Out;

	assign add_kernel2=channel1_Kernel2_Valid_Out & channel2_Kernel2_Valid_Out & channel3_Kernel2_Valid_Out & channel4_Kernel2_Valid_Out & channel5_Kernel2_Valid_Out & channel6_Kernel2_Valid_Out & channel7_Kernel2_Valid_Out & channel8_Kernel2_Valid_Out & channel9_Kernel2_Valid_Out & channel10_Kernel2_Valid_Out & channel11_Kernel2_Valid_Out & channel12_Kernel2_Valid_Out & channel13_Kernel2_Valid_Out & channel14_Kernel2_Valid_Out & channel15_Kernel2_Valid_Out & channel16_Kernel2_Valid_Out & channel17_Kernel2_Valid_Out & channel18_Kernel2_Valid_Out & channel19_Kernel2_Valid_Out & channel20_Kernel2_Valid_Out & channel21_Kernel2_Valid_Out & channel22_Kernel2_Valid_Out & channel23_Kernel2_Valid_Out & channel24_Kernel2_Valid_Out & channel25_Kernel2_Valid_Out & channel26_Kernel2_Valid_Out & channel27_Kernel2_Valid_Out & channel28_Kernel2_Valid_Out & channel29_Kernel2_Valid_Out & channel30_Kernel2_Valid_Out & channel31_Kernel2_Valid_Out & channel32_Kernel2_Valid_Out;

	wire channel1_Kernel3_Valid_Out, channel2_Kernel3_Valid_Out, channel3_Kernel3_Valid_Out, channel4_Kernel3_Valid_Out, channel5_Kernel3_Valid_Out, channel6_Kernel3_Valid_Out, channel7_Kernel3_Valid_Out, channel8_Kernel3_Valid_Out, channel9_Kernel3_Valid_Out, channel10_Kernel3_Valid_Out, channel11_Kernel3_Valid_Out, channel12_Kernel3_Valid_Out, channel13_Kernel3_Valid_Out, channel14_Kernel3_Valid_Out, channel15_Kernel3_Valid_Out, channel16_Kernel3_Valid_Out, channel17_Kernel3_Valid_Out, channel18_Kernel3_Valid_Out, channel19_Kernel3_Valid_Out, channel20_Kernel3_Valid_Out, channel21_Kernel3_Valid_Out, channel22_Kernel3_Valid_Out, channel23_Kernel3_Valid_Out, channel24_Kernel3_Valid_Out, channel25_Kernel3_Valid_Out, channel26_Kernel3_Valid_Out, channel27_Kernel3_Valid_Out, channel28_Kernel3_Valid_Out, channel29_Kernel3_Valid_Out, channel30_Kernel3_Valid_Out, channel31_Kernel3_Valid_Out, channel32_Kernel3_Valid_Out;

	assign add_kernel3=channel1_Kernel3_Valid_Out & channel2_Kernel3_Valid_Out & channel3_Kernel3_Valid_Out & channel4_Kernel3_Valid_Out & channel5_Kernel3_Valid_Out & channel6_Kernel3_Valid_Out & channel7_Kernel3_Valid_Out & channel8_Kernel3_Valid_Out & channel9_Kernel3_Valid_Out & channel10_Kernel3_Valid_Out & channel11_Kernel3_Valid_Out & channel12_Kernel3_Valid_Out & channel13_Kernel3_Valid_Out & channel14_Kernel3_Valid_Out & channel15_Kernel3_Valid_Out & channel16_Kernel3_Valid_Out & channel17_Kernel3_Valid_Out & channel18_Kernel3_Valid_Out & channel19_Kernel3_Valid_Out & channel20_Kernel3_Valid_Out & channel21_Kernel3_Valid_Out & channel22_Kernel3_Valid_Out & channel23_Kernel3_Valid_Out & channel24_Kernel3_Valid_Out & channel25_Kernel3_Valid_Out & channel26_Kernel3_Valid_Out & channel27_Kernel3_Valid_Out & channel28_Kernel3_Valid_Out & channel29_Kernel3_Valid_Out & channel30_Kernel3_Valid_Out & channel31_Kernel3_Valid_Out & channel32_Kernel3_Valid_Out;

	wire channel1_Kernel4_Valid_Out, channel2_Kernel4_Valid_Out, channel3_Kernel4_Valid_Out, channel4_Kernel4_Valid_Out, channel5_Kernel4_Valid_Out, channel6_Kernel4_Valid_Out, channel7_Kernel4_Valid_Out, channel8_Kernel4_Valid_Out, channel9_Kernel4_Valid_Out, channel10_Kernel4_Valid_Out, channel11_Kernel4_Valid_Out, channel12_Kernel4_Valid_Out, channel13_Kernel4_Valid_Out, channel14_Kernel4_Valid_Out, channel15_Kernel4_Valid_Out, channel16_Kernel4_Valid_Out, channel17_Kernel4_Valid_Out, channel18_Kernel4_Valid_Out, channel19_Kernel4_Valid_Out, channel20_Kernel4_Valid_Out, channel21_Kernel4_Valid_Out, channel22_Kernel4_Valid_Out, channel23_Kernel4_Valid_Out, channel24_Kernel4_Valid_Out, channel25_Kernel4_Valid_Out, channel26_Kernel4_Valid_Out, channel27_Kernel4_Valid_Out, channel28_Kernel4_Valid_Out, channel29_Kernel4_Valid_Out, channel30_Kernel4_Valid_Out, channel31_Kernel4_Valid_Out, channel32_Kernel4_Valid_Out;

	assign add_kernel4=channel1_Kernel4_Valid_Out & channel2_Kernel4_Valid_Out & channel3_Kernel4_Valid_Out & channel4_Kernel4_Valid_Out & channel5_Kernel4_Valid_Out & channel6_Kernel4_Valid_Out & channel7_Kernel4_Valid_Out & channel8_Kernel4_Valid_Out & channel9_Kernel4_Valid_Out & channel10_Kernel4_Valid_Out & channel11_Kernel4_Valid_Out & channel12_Kernel4_Valid_Out & channel13_Kernel4_Valid_Out & channel14_Kernel4_Valid_Out & channel15_Kernel4_Valid_Out & channel16_Kernel4_Valid_Out & channel17_Kernel4_Valid_Out & channel18_Kernel4_Valid_Out & channel19_Kernel4_Valid_Out & channel20_Kernel4_Valid_Out & channel21_Kernel4_Valid_Out & channel22_Kernel4_Valid_Out & channel23_Kernel4_Valid_Out & channel24_Kernel4_Valid_Out & channel25_Kernel4_Valid_Out & channel26_Kernel4_Valid_Out & channel27_Kernel4_Valid_Out & channel28_Kernel4_Valid_Out & channel29_Kernel4_Valid_Out & channel30_Kernel4_Valid_Out & channel31_Kernel4_Valid_Out & channel32_Kernel4_Valid_Out;

	wire channel1_Kernel5_Valid_Out, channel2_Kernel5_Valid_Out, channel3_Kernel5_Valid_Out, channel4_Kernel5_Valid_Out, channel5_Kernel5_Valid_Out, channel6_Kernel5_Valid_Out, channel7_Kernel5_Valid_Out, channel8_Kernel5_Valid_Out, channel9_Kernel5_Valid_Out, channel10_Kernel5_Valid_Out, channel11_Kernel5_Valid_Out, channel12_Kernel5_Valid_Out, channel13_Kernel5_Valid_Out, channel14_Kernel5_Valid_Out, channel15_Kernel5_Valid_Out, channel16_Kernel5_Valid_Out, channel17_Kernel5_Valid_Out, channel18_Kernel5_Valid_Out, channel19_Kernel5_Valid_Out, channel20_Kernel5_Valid_Out, channel21_Kernel5_Valid_Out, channel22_Kernel5_Valid_Out, channel23_Kernel5_Valid_Out, channel24_Kernel5_Valid_Out, channel25_Kernel5_Valid_Out, channel26_Kernel5_Valid_Out, channel27_Kernel5_Valid_Out, channel28_Kernel5_Valid_Out, channel29_Kernel5_Valid_Out, channel30_Kernel5_Valid_Out, channel31_Kernel5_Valid_Out, channel32_Kernel5_Valid_Out;

	assign add_kernel5=channel1_Kernel5_Valid_Out & channel2_Kernel5_Valid_Out & channel3_Kernel5_Valid_Out & channel4_Kernel5_Valid_Out & channel5_Kernel5_Valid_Out & channel6_Kernel5_Valid_Out & channel7_Kernel5_Valid_Out & channel8_Kernel5_Valid_Out & channel9_Kernel5_Valid_Out & channel10_Kernel5_Valid_Out & channel11_Kernel5_Valid_Out & channel12_Kernel5_Valid_Out & channel13_Kernel5_Valid_Out & channel14_Kernel5_Valid_Out & channel15_Kernel5_Valid_Out & channel16_Kernel5_Valid_Out & channel17_Kernel5_Valid_Out & channel18_Kernel5_Valid_Out & channel19_Kernel5_Valid_Out & channel20_Kernel5_Valid_Out & channel21_Kernel5_Valid_Out & channel22_Kernel5_Valid_Out & channel23_Kernel5_Valid_Out & channel24_Kernel5_Valid_Out & channel25_Kernel5_Valid_Out & channel26_Kernel5_Valid_Out & channel27_Kernel5_Valid_Out & channel28_Kernel5_Valid_Out & channel29_Kernel5_Valid_Out & channel30_Kernel5_Valid_Out & channel31_Kernel5_Valid_Out & channel32_Kernel5_Valid_Out;

	wire channel1_Kernel6_Valid_Out, channel2_Kernel6_Valid_Out, channel3_Kernel6_Valid_Out, channel4_Kernel6_Valid_Out, channel5_Kernel6_Valid_Out, channel6_Kernel6_Valid_Out, channel7_Kernel6_Valid_Out, channel8_Kernel6_Valid_Out, channel9_Kernel6_Valid_Out, channel10_Kernel6_Valid_Out, channel11_Kernel6_Valid_Out, channel12_Kernel6_Valid_Out, channel13_Kernel6_Valid_Out, channel14_Kernel6_Valid_Out, channel15_Kernel6_Valid_Out, channel16_Kernel6_Valid_Out, channel17_Kernel6_Valid_Out, channel18_Kernel6_Valid_Out, channel19_Kernel6_Valid_Out, channel20_Kernel6_Valid_Out, channel21_Kernel6_Valid_Out, channel22_Kernel6_Valid_Out, channel23_Kernel6_Valid_Out, channel24_Kernel6_Valid_Out, channel25_Kernel6_Valid_Out, channel26_Kernel6_Valid_Out, channel27_Kernel6_Valid_Out, channel28_Kernel6_Valid_Out, channel29_Kernel6_Valid_Out, channel30_Kernel6_Valid_Out, channel31_Kernel6_Valid_Out, channel32_Kernel6_Valid_Out;

	assign add_kernel6=channel1_Kernel6_Valid_Out & channel2_Kernel6_Valid_Out & channel3_Kernel6_Valid_Out & channel4_Kernel6_Valid_Out & channel5_Kernel6_Valid_Out & channel6_Kernel6_Valid_Out & channel7_Kernel6_Valid_Out & channel8_Kernel6_Valid_Out & channel9_Kernel6_Valid_Out & channel10_Kernel6_Valid_Out & channel11_Kernel6_Valid_Out & channel12_Kernel6_Valid_Out & channel13_Kernel6_Valid_Out & channel14_Kernel6_Valid_Out & channel15_Kernel6_Valid_Out & channel16_Kernel6_Valid_Out & channel17_Kernel6_Valid_Out & channel18_Kernel6_Valid_Out & channel19_Kernel6_Valid_Out & channel20_Kernel6_Valid_Out & channel21_Kernel6_Valid_Out & channel22_Kernel6_Valid_Out & channel23_Kernel6_Valid_Out & channel24_Kernel6_Valid_Out & channel25_Kernel6_Valid_Out & channel26_Kernel6_Valid_Out & channel27_Kernel6_Valid_Out & channel28_Kernel6_Valid_Out & channel29_Kernel6_Valid_Out & channel30_Kernel6_Valid_Out & channel31_Kernel6_Valid_Out & channel32_Kernel6_Valid_Out;

	wire channel1_Kernel7_Valid_Out, channel2_Kernel7_Valid_Out, channel3_Kernel7_Valid_Out, channel4_Kernel7_Valid_Out, channel5_Kernel7_Valid_Out, channel6_Kernel7_Valid_Out, channel7_Kernel7_Valid_Out, channel8_Kernel7_Valid_Out, channel9_Kernel7_Valid_Out, channel10_Kernel7_Valid_Out, channel11_Kernel7_Valid_Out, channel12_Kernel7_Valid_Out, channel13_Kernel7_Valid_Out, channel14_Kernel7_Valid_Out, channel15_Kernel7_Valid_Out, channel16_Kernel7_Valid_Out, channel17_Kernel7_Valid_Out, channel18_Kernel7_Valid_Out, channel19_Kernel7_Valid_Out, channel20_Kernel7_Valid_Out, channel21_Kernel7_Valid_Out, channel22_Kernel7_Valid_Out, channel23_Kernel7_Valid_Out, channel24_Kernel7_Valid_Out, channel25_Kernel7_Valid_Out, channel26_Kernel7_Valid_Out, channel27_Kernel7_Valid_Out, channel28_Kernel7_Valid_Out, channel29_Kernel7_Valid_Out, channel30_Kernel7_Valid_Out, channel31_Kernel7_Valid_Out, channel32_Kernel7_Valid_Out;

	assign add_kernel7=channel1_Kernel7_Valid_Out & channel2_Kernel7_Valid_Out & channel3_Kernel7_Valid_Out & channel4_Kernel7_Valid_Out & channel5_Kernel7_Valid_Out & channel6_Kernel7_Valid_Out & channel7_Kernel7_Valid_Out & channel8_Kernel7_Valid_Out & channel9_Kernel7_Valid_Out & channel10_Kernel7_Valid_Out & channel11_Kernel7_Valid_Out & channel12_Kernel7_Valid_Out & channel13_Kernel7_Valid_Out & channel14_Kernel7_Valid_Out & channel15_Kernel7_Valid_Out & channel16_Kernel7_Valid_Out & channel17_Kernel7_Valid_Out & channel18_Kernel7_Valid_Out & channel19_Kernel7_Valid_Out & channel20_Kernel7_Valid_Out & channel21_Kernel7_Valid_Out & channel22_Kernel7_Valid_Out & channel23_Kernel7_Valid_Out & channel24_Kernel7_Valid_Out & channel25_Kernel7_Valid_Out & channel26_Kernel7_Valid_Out & channel27_Kernel7_Valid_Out & channel28_Kernel7_Valid_Out & channel29_Kernel7_Valid_Out & channel30_Kernel7_Valid_Out & channel31_Kernel7_Valid_Out & channel32_Kernel7_Valid_Out;

	wire channel1_Kernel8_Valid_Out, channel2_Kernel8_Valid_Out, channel3_Kernel8_Valid_Out, channel4_Kernel8_Valid_Out, channel5_Kernel8_Valid_Out, channel6_Kernel8_Valid_Out, channel7_Kernel8_Valid_Out, channel8_Kernel8_Valid_Out, channel9_Kernel8_Valid_Out, channel10_Kernel8_Valid_Out, channel11_Kernel8_Valid_Out, channel12_Kernel8_Valid_Out, channel13_Kernel8_Valid_Out, channel14_Kernel8_Valid_Out, channel15_Kernel8_Valid_Out, channel16_Kernel8_Valid_Out, channel17_Kernel8_Valid_Out, channel18_Kernel8_Valid_Out, channel19_Kernel8_Valid_Out, channel20_Kernel8_Valid_Out, channel21_Kernel8_Valid_Out, channel22_Kernel8_Valid_Out, channel23_Kernel8_Valid_Out, channel24_Kernel8_Valid_Out, channel25_Kernel8_Valid_Out, channel26_Kernel8_Valid_Out, channel27_Kernel8_Valid_Out, channel28_Kernel8_Valid_Out, channel29_Kernel8_Valid_Out, channel30_Kernel8_Valid_Out, channel31_Kernel8_Valid_Out, channel32_Kernel8_Valid_Out;

	assign add_kernel8=channel1_Kernel8_Valid_Out & channel2_Kernel8_Valid_Out & channel3_Kernel8_Valid_Out & channel4_Kernel8_Valid_Out & channel5_Kernel8_Valid_Out & channel6_Kernel8_Valid_Out & channel7_Kernel8_Valid_Out & channel8_Kernel8_Valid_Out & channel9_Kernel8_Valid_Out & channel10_Kernel8_Valid_Out & channel11_Kernel8_Valid_Out & channel12_Kernel8_Valid_Out & channel13_Kernel8_Valid_Out & channel14_Kernel8_Valid_Out & channel15_Kernel8_Valid_Out & channel16_Kernel8_Valid_Out & channel17_Kernel8_Valid_Out & channel18_Kernel8_Valid_Out & channel19_Kernel8_Valid_Out & channel20_Kernel8_Valid_Out & channel21_Kernel8_Valid_Out & channel22_Kernel8_Valid_Out & channel23_Kernel8_Valid_Out & channel24_Kernel8_Valid_Out & channel25_Kernel8_Valid_Out & channel26_Kernel8_Valid_Out & channel27_Kernel8_Valid_Out & channel28_Kernel8_Valid_Out & channel29_Kernel8_Valid_Out & channel30_Kernel8_Valid_Out & channel31_Kernel8_Valid_Out & channel32_Kernel8_Valid_Out;

	wire channel1_Kernel9_Valid_Out, channel2_Kernel9_Valid_Out, channel3_Kernel9_Valid_Out, channel4_Kernel9_Valid_Out, channel5_Kernel9_Valid_Out, channel6_Kernel9_Valid_Out, channel7_Kernel9_Valid_Out, channel8_Kernel9_Valid_Out, channel9_Kernel9_Valid_Out, channel10_Kernel9_Valid_Out, channel11_Kernel9_Valid_Out, channel12_Kernel9_Valid_Out, channel13_Kernel9_Valid_Out, channel14_Kernel9_Valid_Out, channel15_Kernel9_Valid_Out, channel16_Kernel9_Valid_Out, channel17_Kernel9_Valid_Out, channel18_Kernel9_Valid_Out, channel19_Kernel9_Valid_Out, channel20_Kernel9_Valid_Out, channel21_Kernel9_Valid_Out, channel22_Kernel9_Valid_Out, channel23_Kernel9_Valid_Out, channel24_Kernel9_Valid_Out, channel25_Kernel9_Valid_Out, channel26_Kernel9_Valid_Out, channel27_Kernel9_Valid_Out, channel28_Kernel9_Valid_Out, channel29_Kernel9_Valid_Out, channel30_Kernel9_Valid_Out, channel31_Kernel9_Valid_Out, channel32_Kernel9_Valid_Out;

	assign add_kernel9=channel1_Kernel9_Valid_Out & channel2_Kernel9_Valid_Out & channel3_Kernel9_Valid_Out & channel4_Kernel9_Valid_Out & channel5_Kernel9_Valid_Out & channel6_Kernel9_Valid_Out & channel7_Kernel9_Valid_Out & channel8_Kernel9_Valid_Out & channel9_Kernel9_Valid_Out & channel10_Kernel9_Valid_Out & channel11_Kernel9_Valid_Out & channel12_Kernel9_Valid_Out & channel13_Kernel9_Valid_Out & channel14_Kernel9_Valid_Out & channel15_Kernel9_Valid_Out & channel16_Kernel9_Valid_Out & channel17_Kernel9_Valid_Out & channel18_Kernel9_Valid_Out & channel19_Kernel9_Valid_Out & channel20_Kernel9_Valid_Out & channel21_Kernel9_Valid_Out & channel22_Kernel9_Valid_Out & channel23_Kernel9_Valid_Out & channel24_Kernel9_Valid_Out & channel25_Kernel9_Valid_Out & channel26_Kernel9_Valid_Out & channel27_Kernel9_Valid_Out & channel28_Kernel9_Valid_Out & channel29_Kernel9_Valid_Out & channel30_Kernel9_Valid_Out & channel31_Kernel9_Valid_Out & channel32_Kernel9_Valid_Out;

	wire channel1_Kernel10_Valid_Out, channel2_Kernel10_Valid_Out, channel3_Kernel10_Valid_Out, channel4_Kernel10_Valid_Out, channel5_Kernel10_Valid_Out, channel6_Kernel10_Valid_Out, channel7_Kernel10_Valid_Out, channel8_Kernel10_Valid_Out, channel9_Kernel10_Valid_Out, channel10_Kernel10_Valid_Out, channel11_Kernel10_Valid_Out, channel12_Kernel10_Valid_Out, channel13_Kernel10_Valid_Out, channel14_Kernel10_Valid_Out, channel15_Kernel10_Valid_Out, channel16_Kernel10_Valid_Out, channel17_Kernel10_Valid_Out, channel18_Kernel10_Valid_Out, channel19_Kernel10_Valid_Out, channel20_Kernel10_Valid_Out, channel21_Kernel10_Valid_Out, channel22_Kernel10_Valid_Out, channel23_Kernel10_Valid_Out, channel24_Kernel10_Valid_Out, channel25_Kernel10_Valid_Out, channel26_Kernel10_Valid_Out, channel27_Kernel10_Valid_Out, channel28_Kernel10_Valid_Out, channel29_Kernel10_Valid_Out, channel30_Kernel10_Valid_Out, channel31_Kernel10_Valid_Out, channel32_Kernel10_Valid_Out;

	assign add_kernel10=channel1_Kernel10_Valid_Out & channel2_Kernel10_Valid_Out & channel3_Kernel10_Valid_Out & channel4_Kernel10_Valid_Out & channel5_Kernel10_Valid_Out & channel6_Kernel10_Valid_Out & channel7_Kernel10_Valid_Out & channel8_Kernel10_Valid_Out & channel9_Kernel10_Valid_Out & channel10_Kernel10_Valid_Out & channel11_Kernel10_Valid_Out & channel12_Kernel10_Valid_Out & channel13_Kernel10_Valid_Out & channel14_Kernel10_Valid_Out & channel15_Kernel10_Valid_Out & channel16_Kernel10_Valid_Out & channel17_Kernel10_Valid_Out & channel18_Kernel10_Valid_Out & channel19_Kernel10_Valid_Out & channel20_Kernel10_Valid_Out & channel21_Kernel10_Valid_Out & channel22_Kernel10_Valid_Out & channel23_Kernel10_Valid_Out & channel24_Kernel10_Valid_Out & channel25_Kernel10_Valid_Out & channel26_Kernel10_Valid_Out & channel27_Kernel10_Valid_Out & channel28_Kernel10_Valid_Out & channel29_Kernel10_Valid_Out & channel30_Kernel10_Valid_Out & channel31_Kernel10_Valid_Out & channel32_Kernel10_Valid_Out;

	wire channel1_Kernel11_Valid_Out, channel2_Kernel11_Valid_Out, channel3_Kernel11_Valid_Out, channel4_Kernel11_Valid_Out, channel5_Kernel11_Valid_Out, channel6_Kernel11_Valid_Out, channel7_Kernel11_Valid_Out, channel8_Kernel11_Valid_Out, channel9_Kernel11_Valid_Out, channel10_Kernel11_Valid_Out, channel11_Kernel11_Valid_Out, channel12_Kernel11_Valid_Out, channel13_Kernel11_Valid_Out, channel14_Kernel11_Valid_Out, channel15_Kernel11_Valid_Out, channel16_Kernel11_Valid_Out, channel17_Kernel11_Valid_Out, channel18_Kernel11_Valid_Out, channel19_Kernel11_Valid_Out, channel20_Kernel11_Valid_Out, channel21_Kernel11_Valid_Out, channel22_Kernel11_Valid_Out, channel23_Kernel11_Valid_Out, channel24_Kernel11_Valid_Out, channel25_Kernel11_Valid_Out, channel26_Kernel11_Valid_Out, channel27_Kernel11_Valid_Out, channel28_Kernel11_Valid_Out, channel29_Kernel11_Valid_Out, channel30_Kernel11_Valid_Out, channel31_Kernel11_Valid_Out, channel32_Kernel11_Valid_Out;

	assign add_kernel11=channel1_Kernel11_Valid_Out & channel2_Kernel11_Valid_Out & channel3_Kernel11_Valid_Out & channel4_Kernel11_Valid_Out & channel5_Kernel11_Valid_Out & channel6_Kernel11_Valid_Out & channel7_Kernel11_Valid_Out & channel8_Kernel11_Valid_Out & channel9_Kernel11_Valid_Out & channel10_Kernel11_Valid_Out & channel11_Kernel11_Valid_Out & channel12_Kernel11_Valid_Out & channel13_Kernel11_Valid_Out & channel14_Kernel11_Valid_Out & channel15_Kernel11_Valid_Out & channel16_Kernel11_Valid_Out & channel17_Kernel11_Valid_Out & channel18_Kernel11_Valid_Out & channel19_Kernel11_Valid_Out & channel20_Kernel11_Valid_Out & channel21_Kernel11_Valid_Out & channel22_Kernel11_Valid_Out & channel23_Kernel11_Valid_Out & channel24_Kernel11_Valid_Out & channel25_Kernel11_Valid_Out & channel26_Kernel11_Valid_Out & channel27_Kernel11_Valid_Out & channel28_Kernel11_Valid_Out & channel29_Kernel11_Valid_Out & channel30_Kernel11_Valid_Out & channel31_Kernel11_Valid_Out & channel32_Kernel11_Valid_Out;

	wire channel1_Kernel12_Valid_Out, channel2_Kernel12_Valid_Out, channel3_Kernel12_Valid_Out, channel4_Kernel12_Valid_Out, channel5_Kernel12_Valid_Out, channel6_Kernel12_Valid_Out, channel7_Kernel12_Valid_Out, channel8_Kernel12_Valid_Out, channel9_Kernel12_Valid_Out, channel10_Kernel12_Valid_Out, channel11_Kernel12_Valid_Out, channel12_Kernel12_Valid_Out, channel13_Kernel12_Valid_Out, channel14_Kernel12_Valid_Out, channel15_Kernel12_Valid_Out, channel16_Kernel12_Valid_Out, channel17_Kernel12_Valid_Out, channel18_Kernel12_Valid_Out, channel19_Kernel12_Valid_Out, channel20_Kernel12_Valid_Out, channel21_Kernel12_Valid_Out, channel22_Kernel12_Valid_Out, channel23_Kernel12_Valid_Out, channel24_Kernel12_Valid_Out, channel25_Kernel12_Valid_Out, channel26_Kernel12_Valid_Out, channel27_Kernel12_Valid_Out, channel28_Kernel12_Valid_Out, channel29_Kernel12_Valid_Out, channel30_Kernel12_Valid_Out, channel31_Kernel12_Valid_Out, channel32_Kernel12_Valid_Out;

	assign add_kernel12=channel1_Kernel12_Valid_Out & channel2_Kernel12_Valid_Out & channel3_Kernel12_Valid_Out & channel4_Kernel12_Valid_Out & channel5_Kernel12_Valid_Out & channel6_Kernel12_Valid_Out & channel7_Kernel12_Valid_Out & channel8_Kernel12_Valid_Out & channel9_Kernel12_Valid_Out & channel10_Kernel12_Valid_Out & channel11_Kernel12_Valid_Out & channel12_Kernel12_Valid_Out & channel13_Kernel12_Valid_Out & channel14_Kernel12_Valid_Out & channel15_Kernel12_Valid_Out & channel16_Kernel12_Valid_Out & channel17_Kernel12_Valid_Out & channel18_Kernel12_Valid_Out & channel19_Kernel12_Valid_Out & channel20_Kernel12_Valid_Out & channel21_Kernel12_Valid_Out & channel22_Kernel12_Valid_Out & channel23_Kernel12_Valid_Out & channel24_Kernel12_Valid_Out & channel25_Kernel12_Valid_Out & channel26_Kernel12_Valid_Out & channel27_Kernel12_Valid_Out & channel28_Kernel12_Valid_Out & channel29_Kernel12_Valid_Out & channel30_Kernel12_Valid_Out & channel31_Kernel12_Valid_Out & channel32_Kernel12_Valid_Out;

	wire channel1_Kernel13_Valid_Out, channel2_Kernel13_Valid_Out, channel3_Kernel13_Valid_Out, channel4_Kernel13_Valid_Out, channel5_Kernel13_Valid_Out, channel6_Kernel13_Valid_Out, channel7_Kernel13_Valid_Out, channel8_Kernel13_Valid_Out, channel9_Kernel13_Valid_Out, channel10_Kernel13_Valid_Out, channel11_Kernel13_Valid_Out, channel12_Kernel13_Valid_Out, channel13_Kernel13_Valid_Out, channel14_Kernel13_Valid_Out, channel15_Kernel13_Valid_Out, channel16_Kernel13_Valid_Out, channel17_Kernel13_Valid_Out, channel18_Kernel13_Valid_Out, channel19_Kernel13_Valid_Out, channel20_Kernel13_Valid_Out, channel21_Kernel13_Valid_Out, channel22_Kernel13_Valid_Out, channel23_Kernel13_Valid_Out, channel24_Kernel13_Valid_Out, channel25_Kernel13_Valid_Out, channel26_Kernel13_Valid_Out, channel27_Kernel13_Valid_Out, channel28_Kernel13_Valid_Out, channel29_Kernel13_Valid_Out, channel30_Kernel13_Valid_Out, channel31_Kernel13_Valid_Out, channel32_Kernel13_Valid_Out;

	assign add_kernel13=channel1_Kernel13_Valid_Out & channel2_Kernel13_Valid_Out & channel3_Kernel13_Valid_Out & channel4_Kernel13_Valid_Out & channel5_Kernel13_Valid_Out & channel6_Kernel13_Valid_Out & channel7_Kernel13_Valid_Out & channel8_Kernel13_Valid_Out & channel9_Kernel13_Valid_Out & channel10_Kernel13_Valid_Out & channel11_Kernel13_Valid_Out & channel12_Kernel13_Valid_Out & channel13_Kernel13_Valid_Out & channel14_Kernel13_Valid_Out & channel15_Kernel13_Valid_Out & channel16_Kernel13_Valid_Out & channel17_Kernel13_Valid_Out & channel18_Kernel13_Valid_Out & channel19_Kernel13_Valid_Out & channel20_Kernel13_Valid_Out & channel21_Kernel13_Valid_Out & channel22_Kernel13_Valid_Out & channel23_Kernel13_Valid_Out & channel24_Kernel13_Valid_Out & channel25_Kernel13_Valid_Out & channel26_Kernel13_Valid_Out & channel27_Kernel13_Valid_Out & channel28_Kernel13_Valid_Out & channel29_Kernel13_Valid_Out & channel30_Kernel13_Valid_Out & channel31_Kernel13_Valid_Out & channel32_Kernel13_Valid_Out;

	wire channel1_Kernel14_Valid_Out, channel2_Kernel14_Valid_Out, channel3_Kernel14_Valid_Out, channel4_Kernel14_Valid_Out, channel5_Kernel14_Valid_Out, channel6_Kernel14_Valid_Out, channel7_Kernel14_Valid_Out, channel8_Kernel14_Valid_Out, channel9_Kernel14_Valid_Out, channel10_Kernel14_Valid_Out, channel11_Kernel14_Valid_Out, channel12_Kernel14_Valid_Out, channel13_Kernel14_Valid_Out, channel14_Kernel14_Valid_Out, channel15_Kernel14_Valid_Out, channel16_Kernel14_Valid_Out, channel17_Kernel14_Valid_Out, channel18_Kernel14_Valid_Out, channel19_Kernel14_Valid_Out, channel20_Kernel14_Valid_Out, channel21_Kernel14_Valid_Out, channel22_Kernel14_Valid_Out, channel23_Kernel14_Valid_Out, channel24_Kernel14_Valid_Out, channel25_Kernel14_Valid_Out, channel26_Kernel14_Valid_Out, channel27_Kernel14_Valid_Out, channel28_Kernel14_Valid_Out, channel29_Kernel14_Valid_Out, channel30_Kernel14_Valid_Out, channel31_Kernel14_Valid_Out, channel32_Kernel14_Valid_Out;

	assign add_kernel14=channel1_Kernel14_Valid_Out & channel2_Kernel14_Valid_Out & channel3_Kernel14_Valid_Out & channel4_Kernel14_Valid_Out & channel5_Kernel14_Valid_Out & channel6_Kernel14_Valid_Out & channel7_Kernel14_Valid_Out & channel8_Kernel14_Valid_Out & channel9_Kernel14_Valid_Out & channel10_Kernel14_Valid_Out & channel11_Kernel14_Valid_Out & channel12_Kernel14_Valid_Out & channel13_Kernel14_Valid_Out & channel14_Kernel14_Valid_Out & channel15_Kernel14_Valid_Out & channel16_Kernel14_Valid_Out & channel17_Kernel14_Valid_Out & channel18_Kernel14_Valid_Out & channel19_Kernel14_Valid_Out & channel20_Kernel14_Valid_Out & channel21_Kernel14_Valid_Out & channel22_Kernel14_Valid_Out & channel23_Kernel14_Valid_Out & channel24_Kernel14_Valid_Out & channel25_Kernel14_Valid_Out & channel26_Kernel14_Valid_Out & channel27_Kernel14_Valid_Out & channel28_Kernel14_Valid_Out & channel29_Kernel14_Valid_Out & channel30_Kernel14_Valid_Out & channel31_Kernel14_Valid_Out & channel32_Kernel14_Valid_Out;

	wire channel1_Kernel15_Valid_Out, channel2_Kernel15_Valid_Out, channel3_Kernel15_Valid_Out, channel4_Kernel15_Valid_Out, channel5_Kernel15_Valid_Out, channel6_Kernel15_Valid_Out, channel7_Kernel15_Valid_Out, channel8_Kernel15_Valid_Out, channel9_Kernel15_Valid_Out, channel10_Kernel15_Valid_Out, channel11_Kernel15_Valid_Out, channel12_Kernel15_Valid_Out, channel13_Kernel15_Valid_Out, channel14_Kernel15_Valid_Out, channel15_Kernel15_Valid_Out, channel16_Kernel15_Valid_Out, channel17_Kernel15_Valid_Out, channel18_Kernel15_Valid_Out, channel19_Kernel15_Valid_Out, channel20_Kernel15_Valid_Out, channel21_Kernel15_Valid_Out, channel22_Kernel15_Valid_Out, channel23_Kernel15_Valid_Out, channel24_Kernel15_Valid_Out, channel25_Kernel15_Valid_Out, channel26_Kernel15_Valid_Out, channel27_Kernel15_Valid_Out, channel28_Kernel15_Valid_Out, channel29_Kernel15_Valid_Out, channel30_Kernel15_Valid_Out, channel31_Kernel15_Valid_Out, channel32_Kernel15_Valid_Out;

	assign add_kernel15=channel1_Kernel15_Valid_Out & channel2_Kernel15_Valid_Out & channel3_Kernel15_Valid_Out & channel4_Kernel15_Valid_Out & channel5_Kernel15_Valid_Out & channel6_Kernel15_Valid_Out & channel7_Kernel15_Valid_Out & channel8_Kernel15_Valid_Out & channel9_Kernel15_Valid_Out & channel10_Kernel15_Valid_Out & channel11_Kernel15_Valid_Out & channel12_Kernel15_Valid_Out & channel13_Kernel15_Valid_Out & channel14_Kernel15_Valid_Out & channel15_Kernel15_Valid_Out & channel16_Kernel15_Valid_Out & channel17_Kernel15_Valid_Out & channel18_Kernel15_Valid_Out & channel19_Kernel15_Valid_Out & channel20_Kernel15_Valid_Out & channel21_Kernel15_Valid_Out & channel22_Kernel15_Valid_Out & channel23_Kernel15_Valid_Out & channel24_Kernel15_Valid_Out & channel25_Kernel15_Valid_Out & channel26_Kernel15_Valid_Out & channel27_Kernel15_Valid_Out & channel28_Kernel15_Valid_Out & channel29_Kernel15_Valid_Out & channel30_Kernel15_Valid_Out & channel31_Kernel15_Valid_Out & channel32_Kernel15_Valid_Out;

	wire channel1_Kernel16_Valid_Out, channel2_Kernel16_Valid_Out, channel3_Kernel16_Valid_Out, channel4_Kernel16_Valid_Out, channel5_Kernel16_Valid_Out, channel6_Kernel16_Valid_Out, channel7_Kernel16_Valid_Out, channel8_Kernel16_Valid_Out, channel9_Kernel16_Valid_Out, channel10_Kernel16_Valid_Out, channel11_Kernel16_Valid_Out, channel12_Kernel16_Valid_Out, channel13_Kernel16_Valid_Out, channel14_Kernel16_Valid_Out, channel15_Kernel16_Valid_Out, channel16_Kernel16_Valid_Out, channel17_Kernel16_Valid_Out, channel18_Kernel16_Valid_Out, channel19_Kernel16_Valid_Out, channel20_Kernel16_Valid_Out, channel21_Kernel16_Valid_Out, channel22_Kernel16_Valid_Out, channel23_Kernel16_Valid_Out, channel24_Kernel16_Valid_Out, channel25_Kernel16_Valid_Out, channel26_Kernel16_Valid_Out, channel27_Kernel16_Valid_Out, channel28_Kernel16_Valid_Out, channel29_Kernel16_Valid_Out, channel30_Kernel16_Valid_Out, channel31_Kernel16_Valid_Out, channel32_Kernel16_Valid_Out;

	assign add_kernel16=channel1_Kernel16_Valid_Out & channel2_Kernel16_Valid_Out & channel3_Kernel16_Valid_Out & channel4_Kernel16_Valid_Out & channel5_Kernel16_Valid_Out & channel6_Kernel16_Valid_Out & channel7_Kernel16_Valid_Out & channel8_Kernel16_Valid_Out & channel9_Kernel16_Valid_Out & channel10_Kernel16_Valid_Out & channel11_Kernel16_Valid_Out & channel12_Kernel16_Valid_Out & channel13_Kernel16_Valid_Out & channel14_Kernel16_Valid_Out & channel15_Kernel16_Valid_Out & channel16_Kernel16_Valid_Out & channel17_Kernel16_Valid_Out & channel18_Kernel16_Valid_Out & channel19_Kernel16_Valid_Out & channel20_Kernel16_Valid_Out & channel21_Kernel16_Valid_Out & channel22_Kernel16_Valid_Out & channel23_Kernel16_Valid_Out & channel24_Kernel16_Valid_Out & channel25_Kernel16_Valid_Out & channel26_Kernel16_Valid_Out & channel27_Kernel16_Valid_Out & channel28_Kernel16_Valid_Out & channel29_Kernel16_Valid_Out & channel30_Kernel16_Valid_Out & channel31_Kernel16_Valid_Out & channel32_Kernel16_Valid_Out;

	wire channel1_Kernel17_Valid_Out, channel2_Kernel17_Valid_Out, channel3_Kernel17_Valid_Out, channel4_Kernel17_Valid_Out, channel5_Kernel17_Valid_Out, channel6_Kernel17_Valid_Out, channel7_Kernel17_Valid_Out, channel8_Kernel17_Valid_Out, channel9_Kernel17_Valid_Out, channel10_Kernel17_Valid_Out, channel11_Kernel17_Valid_Out, channel12_Kernel17_Valid_Out, channel13_Kernel17_Valid_Out, channel14_Kernel17_Valid_Out, channel15_Kernel17_Valid_Out, channel16_Kernel17_Valid_Out, channel17_Kernel17_Valid_Out, channel18_Kernel17_Valid_Out, channel19_Kernel17_Valid_Out, channel20_Kernel17_Valid_Out, channel21_Kernel17_Valid_Out, channel22_Kernel17_Valid_Out, channel23_Kernel17_Valid_Out, channel24_Kernel17_Valid_Out, channel25_Kernel17_Valid_Out, channel26_Kernel17_Valid_Out, channel27_Kernel17_Valid_Out, channel28_Kernel17_Valid_Out, channel29_Kernel17_Valid_Out, channel30_Kernel17_Valid_Out, channel31_Kernel17_Valid_Out, channel32_Kernel17_Valid_Out;

	assign add_kernel17=channel1_Kernel17_Valid_Out & channel2_Kernel17_Valid_Out & channel3_Kernel17_Valid_Out & channel4_Kernel17_Valid_Out & channel5_Kernel17_Valid_Out & channel6_Kernel17_Valid_Out & channel7_Kernel17_Valid_Out & channel8_Kernel17_Valid_Out & channel9_Kernel17_Valid_Out & channel10_Kernel17_Valid_Out & channel11_Kernel17_Valid_Out & channel12_Kernel17_Valid_Out & channel13_Kernel17_Valid_Out & channel14_Kernel17_Valid_Out & channel15_Kernel17_Valid_Out & channel16_Kernel17_Valid_Out & channel17_Kernel17_Valid_Out & channel18_Kernel17_Valid_Out & channel19_Kernel17_Valid_Out & channel20_Kernel17_Valid_Out & channel21_Kernel17_Valid_Out & channel22_Kernel17_Valid_Out & channel23_Kernel17_Valid_Out & channel24_Kernel17_Valid_Out & channel25_Kernel17_Valid_Out & channel26_Kernel17_Valid_Out & channel27_Kernel17_Valid_Out & channel28_Kernel17_Valid_Out & channel29_Kernel17_Valid_Out & channel30_Kernel17_Valid_Out & channel31_Kernel17_Valid_Out & channel32_Kernel17_Valid_Out;

	wire channel1_Kernel18_Valid_Out, channel2_Kernel18_Valid_Out, channel3_Kernel18_Valid_Out, channel4_Kernel18_Valid_Out, channel5_Kernel18_Valid_Out, channel6_Kernel18_Valid_Out, channel7_Kernel18_Valid_Out, channel8_Kernel18_Valid_Out, channel9_Kernel18_Valid_Out, channel10_Kernel18_Valid_Out, channel11_Kernel18_Valid_Out, channel12_Kernel18_Valid_Out, channel13_Kernel18_Valid_Out, channel14_Kernel18_Valid_Out, channel15_Kernel18_Valid_Out, channel16_Kernel18_Valid_Out, channel17_Kernel18_Valid_Out, channel18_Kernel18_Valid_Out, channel19_Kernel18_Valid_Out, channel20_Kernel18_Valid_Out, channel21_Kernel18_Valid_Out, channel22_Kernel18_Valid_Out, channel23_Kernel18_Valid_Out, channel24_Kernel18_Valid_Out, channel25_Kernel18_Valid_Out, channel26_Kernel18_Valid_Out, channel27_Kernel18_Valid_Out, channel28_Kernel18_Valid_Out, channel29_Kernel18_Valid_Out, channel30_Kernel18_Valid_Out, channel31_Kernel18_Valid_Out, channel32_Kernel18_Valid_Out;

	assign add_kernel18=channel1_Kernel18_Valid_Out & channel2_Kernel18_Valid_Out & channel3_Kernel18_Valid_Out & channel4_Kernel18_Valid_Out & channel5_Kernel18_Valid_Out & channel6_Kernel18_Valid_Out & channel7_Kernel18_Valid_Out & channel8_Kernel18_Valid_Out & channel9_Kernel18_Valid_Out & channel10_Kernel18_Valid_Out & channel11_Kernel18_Valid_Out & channel12_Kernel18_Valid_Out & channel13_Kernel18_Valid_Out & channel14_Kernel18_Valid_Out & channel15_Kernel18_Valid_Out & channel16_Kernel18_Valid_Out & channel17_Kernel18_Valid_Out & channel18_Kernel18_Valid_Out & channel19_Kernel18_Valid_Out & channel20_Kernel18_Valid_Out & channel21_Kernel18_Valid_Out & channel22_Kernel18_Valid_Out & channel23_Kernel18_Valid_Out & channel24_Kernel18_Valid_Out & channel25_Kernel18_Valid_Out & channel26_Kernel18_Valid_Out & channel27_Kernel18_Valid_Out & channel28_Kernel18_Valid_Out & channel29_Kernel18_Valid_Out & channel30_Kernel18_Valid_Out & channel31_Kernel18_Valid_Out & channel32_Kernel18_Valid_Out;

	wire channel1_Kernel19_Valid_Out, channel2_Kernel19_Valid_Out, channel3_Kernel19_Valid_Out, channel4_Kernel19_Valid_Out, channel5_Kernel19_Valid_Out, channel6_Kernel19_Valid_Out, channel7_Kernel19_Valid_Out, channel8_Kernel19_Valid_Out, channel9_Kernel19_Valid_Out, channel10_Kernel19_Valid_Out, channel11_Kernel19_Valid_Out, channel12_Kernel19_Valid_Out, channel13_Kernel19_Valid_Out, channel14_Kernel19_Valid_Out, channel15_Kernel19_Valid_Out, channel16_Kernel19_Valid_Out, channel17_Kernel19_Valid_Out, channel18_Kernel19_Valid_Out, channel19_Kernel19_Valid_Out, channel20_Kernel19_Valid_Out, channel21_Kernel19_Valid_Out, channel22_Kernel19_Valid_Out, channel23_Kernel19_Valid_Out, channel24_Kernel19_Valid_Out, channel25_Kernel19_Valid_Out, channel26_Kernel19_Valid_Out, channel27_Kernel19_Valid_Out, channel28_Kernel19_Valid_Out, channel29_Kernel19_Valid_Out, channel30_Kernel19_Valid_Out, channel31_Kernel19_Valid_Out, channel32_Kernel19_Valid_Out;

	assign add_kernel19=channel1_Kernel19_Valid_Out & channel2_Kernel19_Valid_Out & channel3_Kernel19_Valid_Out & channel4_Kernel19_Valid_Out & channel5_Kernel19_Valid_Out & channel6_Kernel19_Valid_Out & channel7_Kernel19_Valid_Out & channel8_Kernel19_Valid_Out & channel9_Kernel19_Valid_Out & channel10_Kernel19_Valid_Out & channel11_Kernel19_Valid_Out & channel12_Kernel19_Valid_Out & channel13_Kernel19_Valid_Out & channel14_Kernel19_Valid_Out & channel15_Kernel19_Valid_Out & channel16_Kernel19_Valid_Out & channel17_Kernel19_Valid_Out & channel18_Kernel19_Valid_Out & channel19_Kernel19_Valid_Out & channel20_Kernel19_Valid_Out & channel21_Kernel19_Valid_Out & channel22_Kernel19_Valid_Out & channel23_Kernel19_Valid_Out & channel24_Kernel19_Valid_Out & channel25_Kernel19_Valid_Out & channel26_Kernel19_Valid_Out & channel27_Kernel19_Valid_Out & channel28_Kernel19_Valid_Out & channel29_Kernel19_Valid_Out & channel30_Kernel19_Valid_Out & channel31_Kernel19_Valid_Out & channel32_Kernel19_Valid_Out;

	wire channel1_Kernel20_Valid_Out, channel2_Kernel20_Valid_Out, channel3_Kernel20_Valid_Out, channel4_Kernel20_Valid_Out, channel5_Kernel20_Valid_Out, channel6_Kernel20_Valid_Out, channel7_Kernel20_Valid_Out, channel8_Kernel20_Valid_Out, channel9_Kernel20_Valid_Out, channel10_Kernel20_Valid_Out, channel11_Kernel20_Valid_Out, channel12_Kernel20_Valid_Out, channel13_Kernel20_Valid_Out, channel14_Kernel20_Valid_Out, channel15_Kernel20_Valid_Out, channel16_Kernel20_Valid_Out, channel17_Kernel20_Valid_Out, channel18_Kernel20_Valid_Out, channel19_Kernel20_Valid_Out, channel20_Kernel20_Valid_Out, channel21_Kernel20_Valid_Out, channel22_Kernel20_Valid_Out, channel23_Kernel20_Valid_Out, channel24_Kernel20_Valid_Out, channel25_Kernel20_Valid_Out, channel26_Kernel20_Valid_Out, channel27_Kernel20_Valid_Out, channel28_Kernel20_Valid_Out, channel29_Kernel20_Valid_Out, channel30_Kernel20_Valid_Out, channel31_Kernel20_Valid_Out, channel32_Kernel20_Valid_Out;

	assign add_kernel20=channel1_Kernel20_Valid_Out & channel2_Kernel20_Valid_Out & channel3_Kernel20_Valid_Out & channel4_Kernel20_Valid_Out & channel5_Kernel20_Valid_Out & channel6_Kernel20_Valid_Out & channel7_Kernel20_Valid_Out & channel8_Kernel20_Valid_Out & channel9_Kernel20_Valid_Out & channel10_Kernel20_Valid_Out & channel11_Kernel20_Valid_Out & channel12_Kernel20_Valid_Out & channel13_Kernel20_Valid_Out & channel14_Kernel20_Valid_Out & channel15_Kernel20_Valid_Out & channel16_Kernel20_Valid_Out & channel17_Kernel20_Valid_Out & channel18_Kernel20_Valid_Out & channel19_Kernel20_Valid_Out & channel20_Kernel20_Valid_Out & channel21_Kernel20_Valid_Out & channel22_Kernel20_Valid_Out & channel23_Kernel20_Valid_Out & channel24_Kernel20_Valid_Out & channel25_Kernel20_Valid_Out & channel26_Kernel20_Valid_Out & channel27_Kernel20_Valid_Out & channel28_Kernel20_Valid_Out & channel29_Kernel20_Valid_Out & channel30_Kernel20_Valid_Out & channel31_Kernel20_Valid_Out & channel32_Kernel20_Valid_Out;

	wire channel1_Kernel21_Valid_Out, channel2_Kernel21_Valid_Out, channel3_Kernel21_Valid_Out, channel4_Kernel21_Valid_Out, channel5_Kernel21_Valid_Out, channel6_Kernel21_Valid_Out, channel7_Kernel21_Valid_Out, channel8_Kernel21_Valid_Out, channel9_Kernel21_Valid_Out, channel10_Kernel21_Valid_Out, channel11_Kernel21_Valid_Out, channel12_Kernel21_Valid_Out, channel13_Kernel21_Valid_Out, channel14_Kernel21_Valid_Out, channel15_Kernel21_Valid_Out, channel16_Kernel21_Valid_Out, channel17_Kernel21_Valid_Out, channel18_Kernel21_Valid_Out, channel19_Kernel21_Valid_Out, channel20_Kernel21_Valid_Out, channel21_Kernel21_Valid_Out, channel22_Kernel21_Valid_Out, channel23_Kernel21_Valid_Out, channel24_Kernel21_Valid_Out, channel25_Kernel21_Valid_Out, channel26_Kernel21_Valid_Out, channel27_Kernel21_Valid_Out, channel28_Kernel21_Valid_Out, channel29_Kernel21_Valid_Out, channel30_Kernel21_Valid_Out, channel31_Kernel21_Valid_Out, channel32_Kernel21_Valid_Out;

	assign add_kernel21=channel1_Kernel21_Valid_Out & channel2_Kernel21_Valid_Out & channel3_Kernel21_Valid_Out & channel4_Kernel21_Valid_Out & channel5_Kernel21_Valid_Out & channel6_Kernel21_Valid_Out & channel7_Kernel21_Valid_Out & channel8_Kernel21_Valid_Out & channel9_Kernel21_Valid_Out & channel10_Kernel21_Valid_Out & channel11_Kernel21_Valid_Out & channel12_Kernel21_Valid_Out & channel13_Kernel21_Valid_Out & channel14_Kernel21_Valid_Out & channel15_Kernel21_Valid_Out & channel16_Kernel21_Valid_Out & channel17_Kernel21_Valid_Out & channel18_Kernel21_Valid_Out & channel19_Kernel21_Valid_Out & channel20_Kernel21_Valid_Out & channel21_Kernel21_Valid_Out & channel22_Kernel21_Valid_Out & channel23_Kernel21_Valid_Out & channel24_Kernel21_Valid_Out & channel25_Kernel21_Valid_Out & channel26_Kernel21_Valid_Out & channel27_Kernel21_Valid_Out & channel28_Kernel21_Valid_Out & channel29_Kernel21_Valid_Out & channel30_Kernel21_Valid_Out & channel31_Kernel21_Valid_Out & channel32_Kernel21_Valid_Out;

	wire channel1_Kernel22_Valid_Out, channel2_Kernel22_Valid_Out, channel3_Kernel22_Valid_Out, channel4_Kernel22_Valid_Out, channel5_Kernel22_Valid_Out, channel6_Kernel22_Valid_Out, channel7_Kernel22_Valid_Out, channel8_Kernel22_Valid_Out, channel9_Kernel22_Valid_Out, channel10_Kernel22_Valid_Out, channel11_Kernel22_Valid_Out, channel12_Kernel22_Valid_Out, channel13_Kernel22_Valid_Out, channel14_Kernel22_Valid_Out, channel15_Kernel22_Valid_Out, channel16_Kernel22_Valid_Out, channel17_Kernel22_Valid_Out, channel18_Kernel22_Valid_Out, channel19_Kernel22_Valid_Out, channel20_Kernel22_Valid_Out, channel21_Kernel22_Valid_Out, channel22_Kernel22_Valid_Out, channel23_Kernel22_Valid_Out, channel24_Kernel22_Valid_Out, channel25_Kernel22_Valid_Out, channel26_Kernel22_Valid_Out, channel27_Kernel22_Valid_Out, channel28_Kernel22_Valid_Out, channel29_Kernel22_Valid_Out, channel30_Kernel22_Valid_Out, channel31_Kernel22_Valid_Out, channel32_Kernel22_Valid_Out;

	assign add_kernel22=channel1_Kernel22_Valid_Out & channel2_Kernel22_Valid_Out & channel3_Kernel22_Valid_Out & channel4_Kernel22_Valid_Out & channel5_Kernel22_Valid_Out & channel6_Kernel22_Valid_Out & channel7_Kernel22_Valid_Out & channel8_Kernel22_Valid_Out & channel9_Kernel22_Valid_Out & channel10_Kernel22_Valid_Out & channel11_Kernel22_Valid_Out & channel12_Kernel22_Valid_Out & channel13_Kernel22_Valid_Out & channel14_Kernel22_Valid_Out & channel15_Kernel22_Valid_Out & channel16_Kernel22_Valid_Out & channel17_Kernel22_Valid_Out & channel18_Kernel22_Valid_Out & channel19_Kernel22_Valid_Out & channel20_Kernel22_Valid_Out & channel21_Kernel22_Valid_Out & channel22_Kernel22_Valid_Out & channel23_Kernel22_Valid_Out & channel24_Kernel22_Valid_Out & channel25_Kernel22_Valid_Out & channel26_Kernel22_Valid_Out & channel27_Kernel22_Valid_Out & channel28_Kernel22_Valid_Out & channel29_Kernel22_Valid_Out & channel30_Kernel22_Valid_Out & channel31_Kernel22_Valid_Out & channel32_Kernel22_Valid_Out;

	wire channel1_Kernel23_Valid_Out, channel2_Kernel23_Valid_Out, channel3_Kernel23_Valid_Out, channel4_Kernel23_Valid_Out, channel5_Kernel23_Valid_Out, channel6_Kernel23_Valid_Out, channel7_Kernel23_Valid_Out, channel8_Kernel23_Valid_Out, channel9_Kernel23_Valid_Out, channel10_Kernel23_Valid_Out, channel11_Kernel23_Valid_Out, channel12_Kernel23_Valid_Out, channel13_Kernel23_Valid_Out, channel14_Kernel23_Valid_Out, channel15_Kernel23_Valid_Out, channel16_Kernel23_Valid_Out, channel17_Kernel23_Valid_Out, channel18_Kernel23_Valid_Out, channel19_Kernel23_Valid_Out, channel20_Kernel23_Valid_Out, channel21_Kernel23_Valid_Out, channel22_Kernel23_Valid_Out, channel23_Kernel23_Valid_Out, channel24_Kernel23_Valid_Out, channel25_Kernel23_Valid_Out, channel26_Kernel23_Valid_Out, channel27_Kernel23_Valid_Out, channel28_Kernel23_Valid_Out, channel29_Kernel23_Valid_Out, channel30_Kernel23_Valid_Out, channel31_Kernel23_Valid_Out, channel32_Kernel23_Valid_Out;

	assign add_kernel23=channel1_Kernel23_Valid_Out & channel2_Kernel23_Valid_Out & channel3_Kernel23_Valid_Out & channel4_Kernel23_Valid_Out & channel5_Kernel23_Valid_Out & channel6_Kernel23_Valid_Out & channel7_Kernel23_Valid_Out & channel8_Kernel23_Valid_Out & channel9_Kernel23_Valid_Out & channel10_Kernel23_Valid_Out & channel11_Kernel23_Valid_Out & channel12_Kernel23_Valid_Out & channel13_Kernel23_Valid_Out & channel14_Kernel23_Valid_Out & channel15_Kernel23_Valid_Out & channel16_Kernel23_Valid_Out & channel17_Kernel23_Valid_Out & channel18_Kernel23_Valid_Out & channel19_Kernel23_Valid_Out & channel20_Kernel23_Valid_Out & channel21_Kernel23_Valid_Out & channel22_Kernel23_Valid_Out & channel23_Kernel23_Valid_Out & channel24_Kernel23_Valid_Out & channel25_Kernel23_Valid_Out & channel26_Kernel23_Valid_Out & channel27_Kernel23_Valid_Out & channel28_Kernel23_Valid_Out & channel29_Kernel23_Valid_Out & channel30_Kernel23_Valid_Out & channel31_Kernel23_Valid_Out & channel32_Kernel23_Valid_Out;

	wire channel1_Kernel24_Valid_Out, channel2_Kernel24_Valid_Out, channel3_Kernel24_Valid_Out, channel4_Kernel24_Valid_Out, channel5_Kernel24_Valid_Out, channel6_Kernel24_Valid_Out, channel7_Kernel24_Valid_Out, channel8_Kernel24_Valid_Out, channel9_Kernel24_Valid_Out, channel10_Kernel24_Valid_Out, channel11_Kernel24_Valid_Out, channel12_Kernel24_Valid_Out, channel13_Kernel24_Valid_Out, channel14_Kernel24_Valid_Out, channel15_Kernel24_Valid_Out, channel16_Kernel24_Valid_Out, channel17_Kernel24_Valid_Out, channel18_Kernel24_Valid_Out, channel19_Kernel24_Valid_Out, channel20_Kernel24_Valid_Out, channel21_Kernel24_Valid_Out, channel22_Kernel24_Valid_Out, channel23_Kernel24_Valid_Out, channel24_Kernel24_Valid_Out, channel25_Kernel24_Valid_Out, channel26_Kernel24_Valid_Out, channel27_Kernel24_Valid_Out, channel28_Kernel24_Valid_Out, channel29_Kernel24_Valid_Out, channel30_Kernel24_Valid_Out, channel31_Kernel24_Valid_Out, channel32_Kernel24_Valid_Out;

	assign add_kernel24=channel1_Kernel24_Valid_Out & channel2_Kernel24_Valid_Out & channel3_Kernel24_Valid_Out & channel4_Kernel24_Valid_Out & channel5_Kernel24_Valid_Out & channel6_Kernel24_Valid_Out & channel7_Kernel24_Valid_Out & channel8_Kernel24_Valid_Out & channel9_Kernel24_Valid_Out & channel10_Kernel24_Valid_Out & channel11_Kernel24_Valid_Out & channel12_Kernel24_Valid_Out & channel13_Kernel24_Valid_Out & channel14_Kernel24_Valid_Out & channel15_Kernel24_Valid_Out & channel16_Kernel24_Valid_Out & channel17_Kernel24_Valid_Out & channel18_Kernel24_Valid_Out & channel19_Kernel24_Valid_Out & channel20_Kernel24_Valid_Out & channel21_Kernel24_Valid_Out & channel22_Kernel24_Valid_Out & channel23_Kernel24_Valid_Out & channel24_Kernel24_Valid_Out & channel25_Kernel24_Valid_Out & channel26_Kernel24_Valid_Out & channel27_Kernel24_Valid_Out & channel28_Kernel24_Valid_Out & channel29_Kernel24_Valid_Out & channel30_Kernel24_Valid_Out & channel31_Kernel24_Valid_Out & channel32_Kernel24_Valid_Out;

	wire channel1_Kernel25_Valid_Out, channel2_Kernel25_Valid_Out, channel3_Kernel25_Valid_Out, channel4_Kernel25_Valid_Out, channel5_Kernel25_Valid_Out, channel6_Kernel25_Valid_Out, channel7_Kernel25_Valid_Out, channel8_Kernel25_Valid_Out, channel9_Kernel25_Valid_Out, channel10_Kernel25_Valid_Out, channel11_Kernel25_Valid_Out, channel12_Kernel25_Valid_Out, channel13_Kernel25_Valid_Out, channel14_Kernel25_Valid_Out, channel15_Kernel25_Valid_Out, channel16_Kernel25_Valid_Out, channel17_Kernel25_Valid_Out, channel18_Kernel25_Valid_Out, channel19_Kernel25_Valid_Out, channel20_Kernel25_Valid_Out, channel21_Kernel25_Valid_Out, channel22_Kernel25_Valid_Out, channel23_Kernel25_Valid_Out, channel24_Kernel25_Valid_Out, channel25_Kernel25_Valid_Out, channel26_Kernel25_Valid_Out, channel27_Kernel25_Valid_Out, channel28_Kernel25_Valid_Out, channel29_Kernel25_Valid_Out, channel30_Kernel25_Valid_Out, channel31_Kernel25_Valid_Out, channel32_Kernel25_Valid_Out;

	assign add_kernel25=channel1_Kernel25_Valid_Out & channel2_Kernel25_Valid_Out & channel3_Kernel25_Valid_Out & channel4_Kernel25_Valid_Out & channel5_Kernel25_Valid_Out & channel6_Kernel25_Valid_Out & channel7_Kernel25_Valid_Out & channel8_Kernel25_Valid_Out & channel9_Kernel25_Valid_Out & channel10_Kernel25_Valid_Out & channel11_Kernel25_Valid_Out & channel12_Kernel25_Valid_Out & channel13_Kernel25_Valid_Out & channel14_Kernel25_Valid_Out & channel15_Kernel25_Valid_Out & channel16_Kernel25_Valid_Out & channel17_Kernel25_Valid_Out & channel18_Kernel25_Valid_Out & channel19_Kernel25_Valid_Out & channel20_Kernel25_Valid_Out & channel21_Kernel25_Valid_Out & channel22_Kernel25_Valid_Out & channel23_Kernel25_Valid_Out & channel24_Kernel25_Valid_Out & channel25_Kernel25_Valid_Out & channel26_Kernel25_Valid_Out & channel27_Kernel25_Valid_Out & channel28_Kernel25_Valid_Out & channel29_Kernel25_Valid_Out & channel30_Kernel25_Valid_Out & channel31_Kernel25_Valid_Out & channel32_Kernel25_Valid_Out;

	wire channel1_Kernel26_Valid_Out, channel2_Kernel26_Valid_Out, channel3_Kernel26_Valid_Out, channel4_Kernel26_Valid_Out, channel5_Kernel26_Valid_Out, channel6_Kernel26_Valid_Out, channel7_Kernel26_Valid_Out, channel8_Kernel26_Valid_Out, channel9_Kernel26_Valid_Out, channel10_Kernel26_Valid_Out, channel11_Kernel26_Valid_Out, channel12_Kernel26_Valid_Out, channel13_Kernel26_Valid_Out, channel14_Kernel26_Valid_Out, channel15_Kernel26_Valid_Out, channel16_Kernel26_Valid_Out, channel17_Kernel26_Valid_Out, channel18_Kernel26_Valid_Out, channel19_Kernel26_Valid_Out, channel20_Kernel26_Valid_Out, channel21_Kernel26_Valid_Out, channel22_Kernel26_Valid_Out, channel23_Kernel26_Valid_Out, channel24_Kernel26_Valid_Out, channel25_Kernel26_Valid_Out, channel26_Kernel26_Valid_Out, channel27_Kernel26_Valid_Out, channel28_Kernel26_Valid_Out, channel29_Kernel26_Valid_Out, channel30_Kernel26_Valid_Out, channel31_Kernel26_Valid_Out, channel32_Kernel26_Valid_Out;

	assign add_kernel26=channel1_Kernel26_Valid_Out & channel2_Kernel26_Valid_Out & channel3_Kernel26_Valid_Out & channel4_Kernel26_Valid_Out & channel5_Kernel26_Valid_Out & channel6_Kernel26_Valid_Out & channel7_Kernel26_Valid_Out & channel8_Kernel26_Valid_Out & channel9_Kernel26_Valid_Out & channel10_Kernel26_Valid_Out & channel11_Kernel26_Valid_Out & channel12_Kernel26_Valid_Out & channel13_Kernel26_Valid_Out & channel14_Kernel26_Valid_Out & channel15_Kernel26_Valid_Out & channel16_Kernel26_Valid_Out & channel17_Kernel26_Valid_Out & channel18_Kernel26_Valid_Out & channel19_Kernel26_Valid_Out & channel20_Kernel26_Valid_Out & channel21_Kernel26_Valid_Out & channel22_Kernel26_Valid_Out & channel23_Kernel26_Valid_Out & channel24_Kernel26_Valid_Out & channel25_Kernel26_Valid_Out & channel26_Kernel26_Valid_Out & channel27_Kernel26_Valid_Out & channel28_Kernel26_Valid_Out & channel29_Kernel26_Valid_Out & channel30_Kernel26_Valid_Out & channel31_Kernel26_Valid_Out & channel32_Kernel26_Valid_Out;

	wire channel1_Kernel27_Valid_Out, channel2_Kernel27_Valid_Out, channel3_Kernel27_Valid_Out, channel4_Kernel27_Valid_Out, channel5_Kernel27_Valid_Out, channel6_Kernel27_Valid_Out, channel7_Kernel27_Valid_Out, channel8_Kernel27_Valid_Out, channel9_Kernel27_Valid_Out, channel10_Kernel27_Valid_Out, channel11_Kernel27_Valid_Out, channel12_Kernel27_Valid_Out, channel13_Kernel27_Valid_Out, channel14_Kernel27_Valid_Out, channel15_Kernel27_Valid_Out, channel16_Kernel27_Valid_Out, channel17_Kernel27_Valid_Out, channel18_Kernel27_Valid_Out, channel19_Kernel27_Valid_Out, channel20_Kernel27_Valid_Out, channel21_Kernel27_Valid_Out, channel22_Kernel27_Valid_Out, channel23_Kernel27_Valid_Out, channel24_Kernel27_Valid_Out, channel25_Kernel27_Valid_Out, channel26_Kernel27_Valid_Out, channel27_Kernel27_Valid_Out, channel28_Kernel27_Valid_Out, channel29_Kernel27_Valid_Out, channel30_Kernel27_Valid_Out, channel31_Kernel27_Valid_Out, channel32_Kernel27_Valid_Out;

	assign add_kernel27=channel1_Kernel27_Valid_Out & channel2_Kernel27_Valid_Out & channel3_Kernel27_Valid_Out & channel4_Kernel27_Valid_Out & channel5_Kernel27_Valid_Out & channel6_Kernel27_Valid_Out & channel7_Kernel27_Valid_Out & channel8_Kernel27_Valid_Out & channel9_Kernel27_Valid_Out & channel10_Kernel27_Valid_Out & channel11_Kernel27_Valid_Out & channel12_Kernel27_Valid_Out & channel13_Kernel27_Valid_Out & channel14_Kernel27_Valid_Out & channel15_Kernel27_Valid_Out & channel16_Kernel27_Valid_Out & channel17_Kernel27_Valid_Out & channel18_Kernel27_Valid_Out & channel19_Kernel27_Valid_Out & channel20_Kernel27_Valid_Out & channel21_Kernel27_Valid_Out & channel22_Kernel27_Valid_Out & channel23_Kernel27_Valid_Out & channel24_Kernel27_Valid_Out & channel25_Kernel27_Valid_Out & channel26_Kernel27_Valid_Out & channel27_Kernel27_Valid_Out & channel28_Kernel27_Valid_Out & channel29_Kernel27_Valid_Out & channel30_Kernel27_Valid_Out & channel31_Kernel27_Valid_Out & channel32_Kernel27_Valid_Out;

	wire channel1_Kernel28_Valid_Out, channel2_Kernel28_Valid_Out, channel3_Kernel28_Valid_Out, channel4_Kernel28_Valid_Out, channel5_Kernel28_Valid_Out, channel6_Kernel28_Valid_Out, channel7_Kernel28_Valid_Out, channel8_Kernel28_Valid_Out, channel9_Kernel28_Valid_Out, channel10_Kernel28_Valid_Out, channel11_Kernel28_Valid_Out, channel12_Kernel28_Valid_Out, channel13_Kernel28_Valid_Out, channel14_Kernel28_Valid_Out, channel15_Kernel28_Valid_Out, channel16_Kernel28_Valid_Out, channel17_Kernel28_Valid_Out, channel18_Kernel28_Valid_Out, channel19_Kernel28_Valid_Out, channel20_Kernel28_Valid_Out, channel21_Kernel28_Valid_Out, channel22_Kernel28_Valid_Out, channel23_Kernel28_Valid_Out, channel24_Kernel28_Valid_Out, channel25_Kernel28_Valid_Out, channel26_Kernel28_Valid_Out, channel27_Kernel28_Valid_Out, channel28_Kernel28_Valid_Out, channel29_Kernel28_Valid_Out, channel30_Kernel28_Valid_Out, channel31_Kernel28_Valid_Out, channel32_Kernel28_Valid_Out;

	assign add_kernel28=channel1_Kernel28_Valid_Out & channel2_Kernel28_Valid_Out & channel3_Kernel28_Valid_Out & channel4_Kernel28_Valid_Out & channel5_Kernel28_Valid_Out & channel6_Kernel28_Valid_Out & channel7_Kernel28_Valid_Out & channel8_Kernel28_Valid_Out & channel9_Kernel28_Valid_Out & channel10_Kernel28_Valid_Out & channel11_Kernel28_Valid_Out & channel12_Kernel28_Valid_Out & channel13_Kernel28_Valid_Out & channel14_Kernel28_Valid_Out & channel15_Kernel28_Valid_Out & channel16_Kernel28_Valid_Out & channel17_Kernel28_Valid_Out & channel18_Kernel28_Valid_Out & channel19_Kernel28_Valid_Out & channel20_Kernel28_Valid_Out & channel21_Kernel28_Valid_Out & channel22_Kernel28_Valid_Out & channel23_Kernel28_Valid_Out & channel24_Kernel28_Valid_Out & channel25_Kernel28_Valid_Out & channel26_Kernel28_Valid_Out & channel27_Kernel28_Valid_Out & channel28_Kernel28_Valid_Out & channel29_Kernel28_Valid_Out & channel30_Kernel28_Valid_Out & channel31_Kernel28_Valid_Out & channel32_Kernel28_Valid_Out;

	wire channel1_Kernel29_Valid_Out, channel2_Kernel29_Valid_Out, channel3_Kernel29_Valid_Out, channel4_Kernel29_Valid_Out, channel5_Kernel29_Valid_Out, channel6_Kernel29_Valid_Out, channel7_Kernel29_Valid_Out, channel8_Kernel29_Valid_Out, channel9_Kernel29_Valid_Out, channel10_Kernel29_Valid_Out, channel11_Kernel29_Valid_Out, channel12_Kernel29_Valid_Out, channel13_Kernel29_Valid_Out, channel14_Kernel29_Valid_Out, channel15_Kernel29_Valid_Out, channel16_Kernel29_Valid_Out, channel17_Kernel29_Valid_Out, channel18_Kernel29_Valid_Out, channel19_Kernel29_Valid_Out, channel20_Kernel29_Valid_Out, channel21_Kernel29_Valid_Out, channel22_Kernel29_Valid_Out, channel23_Kernel29_Valid_Out, channel24_Kernel29_Valid_Out, channel25_Kernel29_Valid_Out, channel26_Kernel29_Valid_Out, channel27_Kernel29_Valid_Out, channel28_Kernel29_Valid_Out, channel29_Kernel29_Valid_Out, channel30_Kernel29_Valid_Out, channel31_Kernel29_Valid_Out, channel32_Kernel29_Valid_Out;

	assign add_kernel29=channel1_Kernel29_Valid_Out & channel2_Kernel29_Valid_Out & channel3_Kernel29_Valid_Out & channel4_Kernel29_Valid_Out & channel5_Kernel29_Valid_Out & channel6_Kernel29_Valid_Out & channel7_Kernel29_Valid_Out & channel8_Kernel29_Valid_Out & channel9_Kernel29_Valid_Out & channel10_Kernel29_Valid_Out & channel11_Kernel29_Valid_Out & channel12_Kernel29_Valid_Out & channel13_Kernel29_Valid_Out & channel14_Kernel29_Valid_Out & channel15_Kernel29_Valid_Out & channel16_Kernel29_Valid_Out & channel17_Kernel29_Valid_Out & channel18_Kernel29_Valid_Out & channel19_Kernel29_Valid_Out & channel20_Kernel29_Valid_Out & channel21_Kernel29_Valid_Out & channel22_Kernel29_Valid_Out & channel23_Kernel29_Valid_Out & channel24_Kernel29_Valid_Out & channel25_Kernel29_Valid_Out & channel26_Kernel29_Valid_Out & channel27_Kernel29_Valid_Out & channel28_Kernel29_Valid_Out & channel29_Kernel29_Valid_Out & channel30_Kernel29_Valid_Out & channel31_Kernel29_Valid_Out & channel32_Kernel29_Valid_Out;

	wire channel1_Kernel30_Valid_Out, channel2_Kernel30_Valid_Out, channel3_Kernel30_Valid_Out, channel4_Kernel30_Valid_Out, channel5_Kernel30_Valid_Out, channel6_Kernel30_Valid_Out, channel7_Kernel30_Valid_Out, channel8_Kernel30_Valid_Out, channel9_Kernel30_Valid_Out, channel10_Kernel30_Valid_Out, channel11_Kernel30_Valid_Out, channel12_Kernel30_Valid_Out, channel13_Kernel30_Valid_Out, channel14_Kernel30_Valid_Out, channel15_Kernel30_Valid_Out, channel16_Kernel30_Valid_Out, channel17_Kernel30_Valid_Out, channel18_Kernel30_Valid_Out, channel19_Kernel30_Valid_Out, channel20_Kernel30_Valid_Out, channel21_Kernel30_Valid_Out, channel22_Kernel30_Valid_Out, channel23_Kernel30_Valid_Out, channel24_Kernel30_Valid_Out, channel25_Kernel30_Valid_Out, channel26_Kernel30_Valid_Out, channel27_Kernel30_Valid_Out, channel28_Kernel30_Valid_Out, channel29_Kernel30_Valid_Out, channel30_Kernel30_Valid_Out, channel31_Kernel30_Valid_Out, channel32_Kernel30_Valid_Out;

	assign add_kernel30=channel1_Kernel30_Valid_Out & channel2_Kernel30_Valid_Out & channel3_Kernel30_Valid_Out & channel4_Kernel30_Valid_Out & channel5_Kernel30_Valid_Out & channel6_Kernel30_Valid_Out & channel7_Kernel30_Valid_Out & channel8_Kernel30_Valid_Out & channel9_Kernel30_Valid_Out & channel10_Kernel30_Valid_Out & channel11_Kernel30_Valid_Out & channel12_Kernel30_Valid_Out & channel13_Kernel30_Valid_Out & channel14_Kernel30_Valid_Out & channel15_Kernel30_Valid_Out & channel16_Kernel30_Valid_Out & channel17_Kernel30_Valid_Out & channel18_Kernel30_Valid_Out & channel19_Kernel30_Valid_Out & channel20_Kernel30_Valid_Out & channel21_Kernel30_Valid_Out & channel22_Kernel30_Valid_Out & channel23_Kernel30_Valid_Out & channel24_Kernel30_Valid_Out & channel25_Kernel30_Valid_Out & channel26_Kernel30_Valid_Out & channel27_Kernel30_Valid_Out & channel28_Kernel30_Valid_Out & channel29_Kernel30_Valid_Out & channel30_Kernel30_Valid_Out & channel31_Kernel30_Valid_Out & channel32_Kernel30_Valid_Out;

	wire channel1_Kernel31_Valid_Out, channel2_Kernel31_Valid_Out, channel3_Kernel31_Valid_Out, channel4_Kernel31_Valid_Out, channel5_Kernel31_Valid_Out, channel6_Kernel31_Valid_Out, channel7_Kernel31_Valid_Out, channel8_Kernel31_Valid_Out, channel9_Kernel31_Valid_Out, channel10_Kernel31_Valid_Out, channel11_Kernel31_Valid_Out, channel12_Kernel31_Valid_Out, channel13_Kernel31_Valid_Out, channel14_Kernel31_Valid_Out, channel15_Kernel31_Valid_Out, channel16_Kernel31_Valid_Out, channel17_Kernel31_Valid_Out, channel18_Kernel31_Valid_Out, channel19_Kernel31_Valid_Out, channel20_Kernel31_Valid_Out, channel21_Kernel31_Valid_Out, channel22_Kernel31_Valid_Out, channel23_Kernel31_Valid_Out, channel24_Kernel31_Valid_Out, channel25_Kernel31_Valid_Out, channel26_Kernel31_Valid_Out, channel27_Kernel31_Valid_Out, channel28_Kernel31_Valid_Out, channel29_Kernel31_Valid_Out, channel30_Kernel31_Valid_Out, channel31_Kernel31_Valid_Out, channel32_Kernel31_Valid_Out;

	assign add_kernel31=channel1_Kernel31_Valid_Out & channel2_Kernel31_Valid_Out & channel3_Kernel31_Valid_Out & channel4_Kernel31_Valid_Out & channel5_Kernel31_Valid_Out & channel6_Kernel31_Valid_Out & channel7_Kernel31_Valid_Out & channel8_Kernel31_Valid_Out & channel9_Kernel31_Valid_Out & channel10_Kernel31_Valid_Out & channel11_Kernel31_Valid_Out & channel12_Kernel31_Valid_Out & channel13_Kernel31_Valid_Out & channel14_Kernel31_Valid_Out & channel15_Kernel31_Valid_Out & channel16_Kernel31_Valid_Out & channel17_Kernel31_Valid_Out & channel18_Kernel31_Valid_Out & channel19_Kernel31_Valid_Out & channel20_Kernel31_Valid_Out & channel21_Kernel31_Valid_Out & channel22_Kernel31_Valid_Out & channel23_Kernel31_Valid_Out & channel24_Kernel31_Valid_Out & channel25_Kernel31_Valid_Out & channel26_Kernel31_Valid_Out & channel27_Kernel31_Valid_Out & channel28_Kernel31_Valid_Out & channel29_Kernel31_Valid_Out & channel30_Kernel31_Valid_Out & channel31_Kernel31_Valid_Out & channel32_Kernel31_Valid_Out;

	wire channel1_Kernel32_Valid_Out, channel2_Kernel32_Valid_Out, channel3_Kernel32_Valid_Out, channel4_Kernel32_Valid_Out, channel5_Kernel32_Valid_Out, channel6_Kernel32_Valid_Out, channel7_Kernel32_Valid_Out, channel8_Kernel32_Valid_Out, channel9_Kernel32_Valid_Out, channel10_Kernel32_Valid_Out, channel11_Kernel32_Valid_Out, channel12_Kernel32_Valid_Out, channel13_Kernel32_Valid_Out, channel14_Kernel32_Valid_Out, channel15_Kernel32_Valid_Out, channel16_Kernel32_Valid_Out, channel17_Kernel32_Valid_Out, channel18_Kernel32_Valid_Out, channel19_Kernel32_Valid_Out, channel20_Kernel32_Valid_Out, channel21_Kernel32_Valid_Out, channel22_Kernel32_Valid_Out, channel23_Kernel32_Valid_Out, channel24_Kernel32_Valid_Out, channel25_Kernel32_Valid_Out, channel26_Kernel32_Valid_Out, channel27_Kernel32_Valid_Out, channel28_Kernel32_Valid_Out, channel29_Kernel32_Valid_Out, channel30_Kernel32_Valid_Out, channel31_Kernel32_Valid_Out, channel32_Kernel32_Valid_Out;

	assign add_kernel32=channel1_Kernel32_Valid_Out & channel2_Kernel32_Valid_Out & channel3_Kernel32_Valid_Out & channel4_Kernel32_Valid_Out & channel5_Kernel32_Valid_Out & channel6_Kernel32_Valid_Out & channel7_Kernel32_Valid_Out & channel8_Kernel32_Valid_Out & channel9_Kernel32_Valid_Out & channel10_Kernel32_Valid_Out & channel11_Kernel32_Valid_Out & channel12_Kernel32_Valid_Out & channel13_Kernel32_Valid_Out & channel14_Kernel32_Valid_Out & channel15_Kernel32_Valid_Out & channel16_Kernel32_Valid_Out & channel17_Kernel32_Valid_Out & channel18_Kernel32_Valid_Out & channel19_Kernel32_Valid_Out & channel20_Kernel32_Valid_Out & channel21_Kernel32_Valid_Out & channel22_Kernel32_Valid_Out & channel23_Kernel32_Valid_Out & channel24_Kernel32_Valid_Out & channel25_Kernel32_Valid_Out & channel26_Kernel32_Valid_Out & channel27_Kernel32_Valid_Out & channel28_Kernel32_Valid_Out & channel29_Kernel32_Valid_Out & channel30_Kernel32_Valid_Out & channel31_Kernel32_Valid_Out & channel32_Kernel32_Valid_Out;

	wire channel1_Kernel33_Valid_Out, channel2_Kernel33_Valid_Out, channel3_Kernel33_Valid_Out, channel4_Kernel33_Valid_Out, channel5_Kernel33_Valid_Out, channel6_Kernel33_Valid_Out, channel7_Kernel33_Valid_Out, channel8_Kernel33_Valid_Out, channel9_Kernel33_Valid_Out, channel10_Kernel33_Valid_Out, channel11_Kernel33_Valid_Out, channel12_Kernel33_Valid_Out, channel13_Kernel33_Valid_Out, channel14_Kernel33_Valid_Out, channel15_Kernel33_Valid_Out, channel16_Kernel33_Valid_Out, channel17_Kernel33_Valid_Out, channel18_Kernel33_Valid_Out, channel19_Kernel33_Valid_Out, channel20_Kernel33_Valid_Out, channel21_Kernel33_Valid_Out, channel22_Kernel33_Valid_Out, channel23_Kernel33_Valid_Out, channel24_Kernel33_Valid_Out, channel25_Kernel33_Valid_Out, channel26_Kernel33_Valid_Out, channel27_Kernel33_Valid_Out, channel28_Kernel33_Valid_Out, channel29_Kernel33_Valid_Out, channel30_Kernel33_Valid_Out, channel31_Kernel33_Valid_Out, channel32_Kernel33_Valid_Out;

	assign add_kernel33=channel1_Kernel33_Valid_Out & channel2_Kernel33_Valid_Out & channel3_Kernel33_Valid_Out & channel4_Kernel33_Valid_Out & channel5_Kernel33_Valid_Out & channel6_Kernel33_Valid_Out & channel7_Kernel33_Valid_Out & channel8_Kernel33_Valid_Out & channel9_Kernel33_Valid_Out & channel10_Kernel33_Valid_Out & channel11_Kernel33_Valid_Out & channel12_Kernel33_Valid_Out & channel13_Kernel33_Valid_Out & channel14_Kernel33_Valid_Out & channel15_Kernel33_Valid_Out & channel16_Kernel33_Valid_Out & channel17_Kernel33_Valid_Out & channel18_Kernel33_Valid_Out & channel19_Kernel33_Valid_Out & channel20_Kernel33_Valid_Out & channel21_Kernel33_Valid_Out & channel22_Kernel33_Valid_Out & channel23_Kernel33_Valid_Out & channel24_Kernel33_Valid_Out & channel25_Kernel33_Valid_Out & channel26_Kernel33_Valid_Out & channel27_Kernel33_Valid_Out & channel28_Kernel33_Valid_Out & channel29_Kernel33_Valid_Out & channel30_Kernel33_Valid_Out & channel31_Kernel33_Valid_Out & channel32_Kernel33_Valid_Out;

	wire channel1_Kernel34_Valid_Out, channel2_Kernel34_Valid_Out, channel3_Kernel34_Valid_Out, channel4_Kernel34_Valid_Out, channel5_Kernel34_Valid_Out, channel6_Kernel34_Valid_Out, channel7_Kernel34_Valid_Out, channel8_Kernel34_Valid_Out, channel9_Kernel34_Valid_Out, channel10_Kernel34_Valid_Out, channel11_Kernel34_Valid_Out, channel12_Kernel34_Valid_Out, channel13_Kernel34_Valid_Out, channel14_Kernel34_Valid_Out, channel15_Kernel34_Valid_Out, channel16_Kernel34_Valid_Out, channel17_Kernel34_Valid_Out, channel18_Kernel34_Valid_Out, channel19_Kernel34_Valid_Out, channel20_Kernel34_Valid_Out, channel21_Kernel34_Valid_Out, channel22_Kernel34_Valid_Out, channel23_Kernel34_Valid_Out, channel24_Kernel34_Valid_Out, channel25_Kernel34_Valid_Out, channel26_Kernel34_Valid_Out, channel27_Kernel34_Valid_Out, channel28_Kernel34_Valid_Out, channel29_Kernel34_Valid_Out, channel30_Kernel34_Valid_Out, channel31_Kernel34_Valid_Out, channel32_Kernel34_Valid_Out;

	assign add_kernel34=channel1_Kernel34_Valid_Out & channel2_Kernel34_Valid_Out & channel3_Kernel34_Valid_Out & channel4_Kernel34_Valid_Out & channel5_Kernel34_Valid_Out & channel6_Kernel34_Valid_Out & channel7_Kernel34_Valid_Out & channel8_Kernel34_Valid_Out & channel9_Kernel34_Valid_Out & channel10_Kernel34_Valid_Out & channel11_Kernel34_Valid_Out & channel12_Kernel34_Valid_Out & channel13_Kernel34_Valid_Out & channel14_Kernel34_Valid_Out & channel15_Kernel34_Valid_Out & channel16_Kernel34_Valid_Out & channel17_Kernel34_Valid_Out & channel18_Kernel34_Valid_Out & channel19_Kernel34_Valid_Out & channel20_Kernel34_Valid_Out & channel21_Kernel34_Valid_Out & channel22_Kernel34_Valid_Out & channel23_Kernel34_Valid_Out & channel24_Kernel34_Valid_Out & channel25_Kernel34_Valid_Out & channel26_Kernel34_Valid_Out & channel27_Kernel34_Valid_Out & channel28_Kernel34_Valid_Out & channel29_Kernel34_Valid_Out & channel30_Kernel34_Valid_Out & channel31_Kernel34_Valid_Out & channel32_Kernel34_Valid_Out;

	wire channel1_Kernel35_Valid_Out, channel2_Kernel35_Valid_Out, channel3_Kernel35_Valid_Out, channel4_Kernel35_Valid_Out, channel5_Kernel35_Valid_Out, channel6_Kernel35_Valid_Out, channel7_Kernel35_Valid_Out, channel8_Kernel35_Valid_Out, channel9_Kernel35_Valid_Out, channel10_Kernel35_Valid_Out, channel11_Kernel35_Valid_Out, channel12_Kernel35_Valid_Out, channel13_Kernel35_Valid_Out, channel14_Kernel35_Valid_Out, channel15_Kernel35_Valid_Out, channel16_Kernel35_Valid_Out, channel17_Kernel35_Valid_Out, channel18_Kernel35_Valid_Out, channel19_Kernel35_Valid_Out, channel20_Kernel35_Valid_Out, channel21_Kernel35_Valid_Out, channel22_Kernel35_Valid_Out, channel23_Kernel35_Valid_Out, channel24_Kernel35_Valid_Out, channel25_Kernel35_Valid_Out, channel26_Kernel35_Valid_Out, channel27_Kernel35_Valid_Out, channel28_Kernel35_Valid_Out, channel29_Kernel35_Valid_Out, channel30_Kernel35_Valid_Out, channel31_Kernel35_Valid_Out, channel32_Kernel35_Valid_Out;

	assign add_kernel35=channel1_Kernel35_Valid_Out & channel2_Kernel35_Valid_Out & channel3_Kernel35_Valid_Out & channel4_Kernel35_Valid_Out & channel5_Kernel35_Valid_Out & channel6_Kernel35_Valid_Out & channel7_Kernel35_Valid_Out & channel8_Kernel35_Valid_Out & channel9_Kernel35_Valid_Out & channel10_Kernel35_Valid_Out & channel11_Kernel35_Valid_Out & channel12_Kernel35_Valid_Out & channel13_Kernel35_Valid_Out & channel14_Kernel35_Valid_Out & channel15_Kernel35_Valid_Out & channel16_Kernel35_Valid_Out & channel17_Kernel35_Valid_Out & channel18_Kernel35_Valid_Out & channel19_Kernel35_Valid_Out & channel20_Kernel35_Valid_Out & channel21_Kernel35_Valid_Out & channel22_Kernel35_Valid_Out & channel23_Kernel35_Valid_Out & channel24_Kernel35_Valid_Out & channel25_Kernel35_Valid_Out & channel26_Kernel35_Valid_Out & channel27_Kernel35_Valid_Out & channel28_Kernel35_Valid_Out & channel29_Kernel35_Valid_Out & channel30_Kernel35_Valid_Out & channel31_Kernel35_Valid_Out & channel32_Kernel35_Valid_Out;

	wire channel1_Kernel36_Valid_Out, channel2_Kernel36_Valid_Out, channel3_Kernel36_Valid_Out, channel4_Kernel36_Valid_Out, channel5_Kernel36_Valid_Out, channel6_Kernel36_Valid_Out, channel7_Kernel36_Valid_Out, channel8_Kernel36_Valid_Out, channel9_Kernel36_Valid_Out, channel10_Kernel36_Valid_Out, channel11_Kernel36_Valid_Out, channel12_Kernel36_Valid_Out, channel13_Kernel36_Valid_Out, channel14_Kernel36_Valid_Out, channel15_Kernel36_Valid_Out, channel16_Kernel36_Valid_Out, channel17_Kernel36_Valid_Out, channel18_Kernel36_Valid_Out, channel19_Kernel36_Valid_Out, channel20_Kernel36_Valid_Out, channel21_Kernel36_Valid_Out, channel22_Kernel36_Valid_Out, channel23_Kernel36_Valid_Out, channel24_Kernel36_Valid_Out, channel25_Kernel36_Valid_Out, channel26_Kernel36_Valid_Out, channel27_Kernel36_Valid_Out, channel28_Kernel36_Valid_Out, channel29_Kernel36_Valid_Out, channel30_Kernel36_Valid_Out, channel31_Kernel36_Valid_Out, channel32_Kernel36_Valid_Out;

	assign add_kernel36=channel1_Kernel36_Valid_Out & channel2_Kernel36_Valid_Out & channel3_Kernel36_Valid_Out & channel4_Kernel36_Valid_Out & channel5_Kernel36_Valid_Out & channel6_Kernel36_Valid_Out & channel7_Kernel36_Valid_Out & channel8_Kernel36_Valid_Out & channel9_Kernel36_Valid_Out & channel10_Kernel36_Valid_Out & channel11_Kernel36_Valid_Out & channel12_Kernel36_Valid_Out & channel13_Kernel36_Valid_Out & channel14_Kernel36_Valid_Out & channel15_Kernel36_Valid_Out & channel16_Kernel36_Valid_Out & channel17_Kernel36_Valid_Out & channel18_Kernel36_Valid_Out & channel19_Kernel36_Valid_Out & channel20_Kernel36_Valid_Out & channel21_Kernel36_Valid_Out & channel22_Kernel36_Valid_Out & channel23_Kernel36_Valid_Out & channel24_Kernel36_Valid_Out & channel25_Kernel36_Valid_Out & channel26_Kernel36_Valid_Out & channel27_Kernel36_Valid_Out & channel28_Kernel36_Valid_Out & channel29_Kernel36_Valid_Out & channel30_Kernel36_Valid_Out & channel31_Kernel36_Valid_Out & channel32_Kernel36_Valid_Out;

	wire channel1_Kernel37_Valid_Out, channel2_Kernel37_Valid_Out, channel3_Kernel37_Valid_Out, channel4_Kernel37_Valid_Out, channel5_Kernel37_Valid_Out, channel6_Kernel37_Valid_Out, channel7_Kernel37_Valid_Out, channel8_Kernel37_Valid_Out, channel9_Kernel37_Valid_Out, channel10_Kernel37_Valid_Out, channel11_Kernel37_Valid_Out, channel12_Kernel37_Valid_Out, channel13_Kernel37_Valid_Out, channel14_Kernel37_Valid_Out, channel15_Kernel37_Valid_Out, channel16_Kernel37_Valid_Out, channel17_Kernel37_Valid_Out, channel18_Kernel37_Valid_Out, channel19_Kernel37_Valid_Out, channel20_Kernel37_Valid_Out, channel21_Kernel37_Valid_Out, channel22_Kernel37_Valid_Out, channel23_Kernel37_Valid_Out, channel24_Kernel37_Valid_Out, channel25_Kernel37_Valid_Out, channel26_Kernel37_Valid_Out, channel27_Kernel37_Valid_Out, channel28_Kernel37_Valid_Out, channel29_Kernel37_Valid_Out, channel30_Kernel37_Valid_Out, channel31_Kernel37_Valid_Out, channel32_Kernel37_Valid_Out;

	assign add_kernel37=channel1_Kernel37_Valid_Out & channel2_Kernel37_Valid_Out & channel3_Kernel37_Valid_Out & channel4_Kernel37_Valid_Out & channel5_Kernel37_Valid_Out & channel6_Kernel37_Valid_Out & channel7_Kernel37_Valid_Out & channel8_Kernel37_Valid_Out & channel9_Kernel37_Valid_Out & channel10_Kernel37_Valid_Out & channel11_Kernel37_Valid_Out & channel12_Kernel37_Valid_Out & channel13_Kernel37_Valid_Out & channel14_Kernel37_Valid_Out & channel15_Kernel37_Valid_Out & channel16_Kernel37_Valid_Out & channel17_Kernel37_Valid_Out & channel18_Kernel37_Valid_Out & channel19_Kernel37_Valid_Out & channel20_Kernel37_Valid_Out & channel21_Kernel37_Valid_Out & channel22_Kernel37_Valid_Out & channel23_Kernel37_Valid_Out & channel24_Kernel37_Valid_Out & channel25_Kernel37_Valid_Out & channel26_Kernel37_Valid_Out & channel27_Kernel37_Valid_Out & channel28_Kernel37_Valid_Out & channel29_Kernel37_Valid_Out & channel30_Kernel37_Valid_Out & channel31_Kernel37_Valid_Out & channel32_Kernel37_Valid_Out;

	wire channel1_Kernel38_Valid_Out, channel2_Kernel38_Valid_Out, channel3_Kernel38_Valid_Out, channel4_Kernel38_Valid_Out, channel5_Kernel38_Valid_Out, channel6_Kernel38_Valid_Out, channel7_Kernel38_Valid_Out, channel8_Kernel38_Valid_Out, channel9_Kernel38_Valid_Out, channel10_Kernel38_Valid_Out, channel11_Kernel38_Valid_Out, channel12_Kernel38_Valid_Out, channel13_Kernel38_Valid_Out, channel14_Kernel38_Valid_Out, channel15_Kernel38_Valid_Out, channel16_Kernel38_Valid_Out, channel17_Kernel38_Valid_Out, channel18_Kernel38_Valid_Out, channel19_Kernel38_Valid_Out, channel20_Kernel38_Valid_Out, channel21_Kernel38_Valid_Out, channel22_Kernel38_Valid_Out, channel23_Kernel38_Valid_Out, channel24_Kernel38_Valid_Out, channel25_Kernel38_Valid_Out, channel26_Kernel38_Valid_Out, channel27_Kernel38_Valid_Out, channel28_Kernel38_Valid_Out, channel29_Kernel38_Valid_Out, channel30_Kernel38_Valid_Out, channel31_Kernel38_Valid_Out, channel32_Kernel38_Valid_Out;

	assign add_kernel38=channel1_Kernel38_Valid_Out & channel2_Kernel38_Valid_Out & channel3_Kernel38_Valid_Out & channel4_Kernel38_Valid_Out & channel5_Kernel38_Valid_Out & channel6_Kernel38_Valid_Out & channel7_Kernel38_Valid_Out & channel8_Kernel38_Valid_Out & channel9_Kernel38_Valid_Out & channel10_Kernel38_Valid_Out & channel11_Kernel38_Valid_Out & channel12_Kernel38_Valid_Out & channel13_Kernel38_Valid_Out & channel14_Kernel38_Valid_Out & channel15_Kernel38_Valid_Out & channel16_Kernel38_Valid_Out & channel17_Kernel38_Valid_Out & channel18_Kernel38_Valid_Out & channel19_Kernel38_Valid_Out & channel20_Kernel38_Valid_Out & channel21_Kernel38_Valid_Out & channel22_Kernel38_Valid_Out & channel23_Kernel38_Valid_Out & channel24_Kernel38_Valid_Out & channel25_Kernel38_Valid_Out & channel26_Kernel38_Valid_Out & channel27_Kernel38_Valid_Out & channel28_Kernel38_Valid_Out & channel29_Kernel38_Valid_Out & channel30_Kernel38_Valid_Out & channel31_Kernel38_Valid_Out & channel32_Kernel38_Valid_Out;

	wire channel1_Kernel39_Valid_Out, channel2_Kernel39_Valid_Out, channel3_Kernel39_Valid_Out, channel4_Kernel39_Valid_Out, channel5_Kernel39_Valid_Out, channel6_Kernel39_Valid_Out, channel7_Kernel39_Valid_Out, channel8_Kernel39_Valid_Out, channel9_Kernel39_Valid_Out, channel10_Kernel39_Valid_Out, channel11_Kernel39_Valid_Out, channel12_Kernel39_Valid_Out, channel13_Kernel39_Valid_Out, channel14_Kernel39_Valid_Out, channel15_Kernel39_Valid_Out, channel16_Kernel39_Valid_Out, channel17_Kernel39_Valid_Out, channel18_Kernel39_Valid_Out, channel19_Kernel39_Valid_Out, channel20_Kernel39_Valid_Out, channel21_Kernel39_Valid_Out, channel22_Kernel39_Valid_Out, channel23_Kernel39_Valid_Out, channel24_Kernel39_Valid_Out, channel25_Kernel39_Valid_Out, channel26_Kernel39_Valid_Out, channel27_Kernel39_Valid_Out, channel28_Kernel39_Valid_Out, channel29_Kernel39_Valid_Out, channel30_Kernel39_Valid_Out, channel31_Kernel39_Valid_Out, channel32_Kernel39_Valid_Out;

	assign add_kernel39=channel1_Kernel39_Valid_Out & channel2_Kernel39_Valid_Out & channel3_Kernel39_Valid_Out & channel4_Kernel39_Valid_Out & channel5_Kernel39_Valid_Out & channel6_Kernel39_Valid_Out & channel7_Kernel39_Valid_Out & channel8_Kernel39_Valid_Out & channel9_Kernel39_Valid_Out & channel10_Kernel39_Valid_Out & channel11_Kernel39_Valid_Out & channel12_Kernel39_Valid_Out & channel13_Kernel39_Valid_Out & channel14_Kernel39_Valid_Out & channel15_Kernel39_Valid_Out & channel16_Kernel39_Valid_Out & channel17_Kernel39_Valid_Out & channel18_Kernel39_Valid_Out & channel19_Kernel39_Valid_Out & channel20_Kernel39_Valid_Out & channel21_Kernel39_Valid_Out & channel22_Kernel39_Valid_Out & channel23_Kernel39_Valid_Out & channel24_Kernel39_Valid_Out & channel25_Kernel39_Valid_Out & channel26_Kernel39_Valid_Out & channel27_Kernel39_Valid_Out & channel28_Kernel39_Valid_Out & channel29_Kernel39_Valid_Out & channel30_Kernel39_Valid_Out & channel31_Kernel39_Valid_Out & channel32_Kernel39_Valid_Out;

	wire channel1_Kernel40_Valid_Out, channel2_Kernel40_Valid_Out, channel3_Kernel40_Valid_Out, channel4_Kernel40_Valid_Out, channel5_Kernel40_Valid_Out, channel6_Kernel40_Valid_Out, channel7_Kernel40_Valid_Out, channel8_Kernel40_Valid_Out, channel9_Kernel40_Valid_Out, channel10_Kernel40_Valid_Out, channel11_Kernel40_Valid_Out, channel12_Kernel40_Valid_Out, channel13_Kernel40_Valid_Out, channel14_Kernel40_Valid_Out, channel15_Kernel40_Valid_Out, channel16_Kernel40_Valid_Out, channel17_Kernel40_Valid_Out, channel18_Kernel40_Valid_Out, channel19_Kernel40_Valid_Out, channel20_Kernel40_Valid_Out, channel21_Kernel40_Valid_Out, channel22_Kernel40_Valid_Out, channel23_Kernel40_Valid_Out, channel24_Kernel40_Valid_Out, channel25_Kernel40_Valid_Out, channel26_Kernel40_Valid_Out, channel27_Kernel40_Valid_Out, channel28_Kernel40_Valid_Out, channel29_Kernel40_Valid_Out, channel30_Kernel40_Valid_Out, channel31_Kernel40_Valid_Out, channel32_Kernel40_Valid_Out;

	assign add_kernel40=channel1_Kernel40_Valid_Out & channel2_Kernel40_Valid_Out & channel3_Kernel40_Valid_Out & channel4_Kernel40_Valid_Out & channel5_Kernel40_Valid_Out & channel6_Kernel40_Valid_Out & channel7_Kernel40_Valid_Out & channel8_Kernel40_Valid_Out & channel9_Kernel40_Valid_Out & channel10_Kernel40_Valid_Out & channel11_Kernel40_Valid_Out & channel12_Kernel40_Valid_Out & channel13_Kernel40_Valid_Out & channel14_Kernel40_Valid_Out & channel15_Kernel40_Valid_Out & channel16_Kernel40_Valid_Out & channel17_Kernel40_Valid_Out & channel18_Kernel40_Valid_Out & channel19_Kernel40_Valid_Out & channel20_Kernel40_Valid_Out & channel21_Kernel40_Valid_Out & channel22_Kernel40_Valid_Out & channel23_Kernel40_Valid_Out & channel24_Kernel40_Valid_Out & channel25_Kernel40_Valid_Out & channel26_Kernel40_Valid_Out & channel27_Kernel40_Valid_Out & channel28_Kernel40_Valid_Out & channel29_Kernel40_Valid_Out & channel30_Kernel40_Valid_Out & channel31_Kernel40_Valid_Out & channel32_Kernel40_Valid_Out;

	wire channel1_Kernel41_Valid_Out, channel2_Kernel41_Valid_Out, channel3_Kernel41_Valid_Out, channel4_Kernel41_Valid_Out, channel5_Kernel41_Valid_Out, channel6_Kernel41_Valid_Out, channel7_Kernel41_Valid_Out, channel8_Kernel41_Valid_Out, channel9_Kernel41_Valid_Out, channel10_Kernel41_Valid_Out, channel11_Kernel41_Valid_Out, channel12_Kernel41_Valid_Out, channel13_Kernel41_Valid_Out, channel14_Kernel41_Valid_Out, channel15_Kernel41_Valid_Out, channel16_Kernel41_Valid_Out, channel17_Kernel41_Valid_Out, channel18_Kernel41_Valid_Out, channel19_Kernel41_Valid_Out, channel20_Kernel41_Valid_Out, channel21_Kernel41_Valid_Out, channel22_Kernel41_Valid_Out, channel23_Kernel41_Valid_Out, channel24_Kernel41_Valid_Out, channel25_Kernel41_Valid_Out, channel26_Kernel41_Valid_Out, channel27_Kernel41_Valid_Out, channel28_Kernel41_Valid_Out, channel29_Kernel41_Valid_Out, channel30_Kernel41_Valid_Out, channel31_Kernel41_Valid_Out, channel32_Kernel41_Valid_Out;

	assign add_kernel41=channel1_Kernel41_Valid_Out & channel2_Kernel41_Valid_Out & channel3_Kernel41_Valid_Out & channel4_Kernel41_Valid_Out & channel5_Kernel41_Valid_Out & channel6_Kernel41_Valid_Out & channel7_Kernel41_Valid_Out & channel8_Kernel41_Valid_Out & channel9_Kernel41_Valid_Out & channel10_Kernel41_Valid_Out & channel11_Kernel41_Valid_Out & channel12_Kernel41_Valid_Out & channel13_Kernel41_Valid_Out & channel14_Kernel41_Valid_Out & channel15_Kernel41_Valid_Out & channel16_Kernel41_Valid_Out & channel17_Kernel41_Valid_Out & channel18_Kernel41_Valid_Out & channel19_Kernel41_Valid_Out & channel20_Kernel41_Valid_Out & channel21_Kernel41_Valid_Out & channel22_Kernel41_Valid_Out & channel23_Kernel41_Valid_Out & channel24_Kernel41_Valid_Out & channel25_Kernel41_Valid_Out & channel26_Kernel41_Valid_Out & channel27_Kernel41_Valid_Out & channel28_Kernel41_Valid_Out & channel29_Kernel41_Valid_Out & channel30_Kernel41_Valid_Out & channel31_Kernel41_Valid_Out & channel32_Kernel41_Valid_Out;

	wire channel1_Kernel42_Valid_Out, channel2_Kernel42_Valid_Out, channel3_Kernel42_Valid_Out, channel4_Kernel42_Valid_Out, channel5_Kernel42_Valid_Out, channel6_Kernel42_Valid_Out, channel7_Kernel42_Valid_Out, channel8_Kernel42_Valid_Out, channel9_Kernel42_Valid_Out, channel10_Kernel42_Valid_Out, channel11_Kernel42_Valid_Out, channel12_Kernel42_Valid_Out, channel13_Kernel42_Valid_Out, channel14_Kernel42_Valid_Out, channel15_Kernel42_Valid_Out, channel16_Kernel42_Valid_Out, channel17_Kernel42_Valid_Out, channel18_Kernel42_Valid_Out, channel19_Kernel42_Valid_Out, channel20_Kernel42_Valid_Out, channel21_Kernel42_Valid_Out, channel22_Kernel42_Valid_Out, channel23_Kernel42_Valid_Out, channel24_Kernel42_Valid_Out, channel25_Kernel42_Valid_Out, channel26_Kernel42_Valid_Out, channel27_Kernel42_Valid_Out, channel28_Kernel42_Valid_Out, channel29_Kernel42_Valid_Out, channel30_Kernel42_Valid_Out, channel31_Kernel42_Valid_Out, channel32_Kernel42_Valid_Out;

	assign add_kernel42=channel1_Kernel42_Valid_Out & channel2_Kernel42_Valid_Out & channel3_Kernel42_Valid_Out & channel4_Kernel42_Valid_Out & channel5_Kernel42_Valid_Out & channel6_Kernel42_Valid_Out & channel7_Kernel42_Valid_Out & channel8_Kernel42_Valid_Out & channel9_Kernel42_Valid_Out & channel10_Kernel42_Valid_Out & channel11_Kernel42_Valid_Out & channel12_Kernel42_Valid_Out & channel13_Kernel42_Valid_Out & channel14_Kernel42_Valid_Out & channel15_Kernel42_Valid_Out & channel16_Kernel42_Valid_Out & channel17_Kernel42_Valid_Out & channel18_Kernel42_Valid_Out & channel19_Kernel42_Valid_Out & channel20_Kernel42_Valid_Out & channel21_Kernel42_Valid_Out & channel22_Kernel42_Valid_Out & channel23_Kernel42_Valid_Out & channel24_Kernel42_Valid_Out & channel25_Kernel42_Valid_Out & channel26_Kernel42_Valid_Out & channel27_Kernel42_Valid_Out & channel28_Kernel42_Valid_Out & channel29_Kernel42_Valid_Out & channel30_Kernel42_Valid_Out & channel31_Kernel42_Valid_Out & channel32_Kernel42_Valid_Out;

	wire channel1_Kernel43_Valid_Out, channel2_Kernel43_Valid_Out, channel3_Kernel43_Valid_Out, channel4_Kernel43_Valid_Out, channel5_Kernel43_Valid_Out, channel6_Kernel43_Valid_Out, channel7_Kernel43_Valid_Out, channel8_Kernel43_Valid_Out, channel9_Kernel43_Valid_Out, channel10_Kernel43_Valid_Out, channel11_Kernel43_Valid_Out, channel12_Kernel43_Valid_Out, channel13_Kernel43_Valid_Out, channel14_Kernel43_Valid_Out, channel15_Kernel43_Valid_Out, channel16_Kernel43_Valid_Out, channel17_Kernel43_Valid_Out, channel18_Kernel43_Valid_Out, channel19_Kernel43_Valid_Out, channel20_Kernel43_Valid_Out, channel21_Kernel43_Valid_Out, channel22_Kernel43_Valid_Out, channel23_Kernel43_Valid_Out, channel24_Kernel43_Valid_Out, channel25_Kernel43_Valid_Out, channel26_Kernel43_Valid_Out, channel27_Kernel43_Valid_Out, channel28_Kernel43_Valid_Out, channel29_Kernel43_Valid_Out, channel30_Kernel43_Valid_Out, channel31_Kernel43_Valid_Out, channel32_Kernel43_Valid_Out;

	assign add_kernel43=channel1_Kernel43_Valid_Out & channel2_Kernel43_Valid_Out & channel3_Kernel43_Valid_Out & channel4_Kernel43_Valid_Out & channel5_Kernel43_Valid_Out & channel6_Kernel43_Valid_Out & channel7_Kernel43_Valid_Out & channel8_Kernel43_Valid_Out & channel9_Kernel43_Valid_Out & channel10_Kernel43_Valid_Out & channel11_Kernel43_Valid_Out & channel12_Kernel43_Valid_Out & channel13_Kernel43_Valid_Out & channel14_Kernel43_Valid_Out & channel15_Kernel43_Valid_Out & channel16_Kernel43_Valid_Out & channel17_Kernel43_Valid_Out & channel18_Kernel43_Valid_Out & channel19_Kernel43_Valid_Out & channel20_Kernel43_Valid_Out & channel21_Kernel43_Valid_Out & channel22_Kernel43_Valid_Out & channel23_Kernel43_Valid_Out & channel24_Kernel43_Valid_Out & channel25_Kernel43_Valid_Out & channel26_Kernel43_Valid_Out & channel27_Kernel43_Valid_Out & channel28_Kernel43_Valid_Out & channel29_Kernel43_Valid_Out & channel30_Kernel43_Valid_Out & channel31_Kernel43_Valid_Out & channel32_Kernel43_Valid_Out;

	wire channel1_Kernel44_Valid_Out, channel2_Kernel44_Valid_Out, channel3_Kernel44_Valid_Out, channel4_Kernel44_Valid_Out, channel5_Kernel44_Valid_Out, channel6_Kernel44_Valid_Out, channel7_Kernel44_Valid_Out, channel8_Kernel44_Valid_Out, channel9_Kernel44_Valid_Out, channel10_Kernel44_Valid_Out, channel11_Kernel44_Valid_Out, channel12_Kernel44_Valid_Out, channel13_Kernel44_Valid_Out, channel14_Kernel44_Valid_Out, channel15_Kernel44_Valid_Out, channel16_Kernel44_Valid_Out, channel17_Kernel44_Valid_Out, channel18_Kernel44_Valid_Out, channel19_Kernel44_Valid_Out, channel20_Kernel44_Valid_Out, channel21_Kernel44_Valid_Out, channel22_Kernel44_Valid_Out, channel23_Kernel44_Valid_Out, channel24_Kernel44_Valid_Out, channel25_Kernel44_Valid_Out, channel26_Kernel44_Valid_Out, channel27_Kernel44_Valid_Out, channel28_Kernel44_Valid_Out, channel29_Kernel44_Valid_Out, channel30_Kernel44_Valid_Out, channel31_Kernel44_Valid_Out, channel32_Kernel44_Valid_Out;

	assign add_kernel44=channel1_Kernel44_Valid_Out & channel2_Kernel44_Valid_Out & channel3_Kernel44_Valid_Out & channel4_Kernel44_Valid_Out & channel5_Kernel44_Valid_Out & channel6_Kernel44_Valid_Out & channel7_Kernel44_Valid_Out & channel8_Kernel44_Valid_Out & channel9_Kernel44_Valid_Out & channel10_Kernel44_Valid_Out & channel11_Kernel44_Valid_Out & channel12_Kernel44_Valid_Out & channel13_Kernel44_Valid_Out & channel14_Kernel44_Valid_Out & channel15_Kernel44_Valid_Out & channel16_Kernel44_Valid_Out & channel17_Kernel44_Valid_Out & channel18_Kernel44_Valid_Out & channel19_Kernel44_Valid_Out & channel20_Kernel44_Valid_Out & channel21_Kernel44_Valid_Out & channel22_Kernel44_Valid_Out & channel23_Kernel44_Valid_Out & channel24_Kernel44_Valid_Out & channel25_Kernel44_Valid_Out & channel26_Kernel44_Valid_Out & channel27_Kernel44_Valid_Out & channel28_Kernel44_Valid_Out & channel29_Kernel44_Valid_Out & channel30_Kernel44_Valid_Out & channel31_Kernel44_Valid_Out & channel32_Kernel44_Valid_Out;

	wire channel1_Kernel45_Valid_Out, channel2_Kernel45_Valid_Out, channel3_Kernel45_Valid_Out, channel4_Kernel45_Valid_Out, channel5_Kernel45_Valid_Out, channel6_Kernel45_Valid_Out, channel7_Kernel45_Valid_Out, channel8_Kernel45_Valid_Out, channel9_Kernel45_Valid_Out, channel10_Kernel45_Valid_Out, channel11_Kernel45_Valid_Out, channel12_Kernel45_Valid_Out, channel13_Kernel45_Valid_Out, channel14_Kernel45_Valid_Out, channel15_Kernel45_Valid_Out, channel16_Kernel45_Valid_Out, channel17_Kernel45_Valid_Out, channel18_Kernel45_Valid_Out, channel19_Kernel45_Valid_Out, channel20_Kernel45_Valid_Out, channel21_Kernel45_Valid_Out, channel22_Kernel45_Valid_Out, channel23_Kernel45_Valid_Out, channel24_Kernel45_Valid_Out, channel25_Kernel45_Valid_Out, channel26_Kernel45_Valid_Out, channel27_Kernel45_Valid_Out, channel28_Kernel45_Valid_Out, channel29_Kernel45_Valid_Out, channel30_Kernel45_Valid_Out, channel31_Kernel45_Valid_Out, channel32_Kernel45_Valid_Out;

	assign add_kernel45=channel1_Kernel45_Valid_Out & channel2_Kernel45_Valid_Out & channel3_Kernel45_Valid_Out & channel4_Kernel45_Valid_Out & channel5_Kernel45_Valid_Out & channel6_Kernel45_Valid_Out & channel7_Kernel45_Valid_Out & channel8_Kernel45_Valid_Out & channel9_Kernel45_Valid_Out & channel10_Kernel45_Valid_Out & channel11_Kernel45_Valid_Out & channel12_Kernel45_Valid_Out & channel13_Kernel45_Valid_Out & channel14_Kernel45_Valid_Out & channel15_Kernel45_Valid_Out & channel16_Kernel45_Valid_Out & channel17_Kernel45_Valid_Out & channel18_Kernel45_Valid_Out & channel19_Kernel45_Valid_Out & channel20_Kernel45_Valid_Out & channel21_Kernel45_Valid_Out & channel22_Kernel45_Valid_Out & channel23_Kernel45_Valid_Out & channel24_Kernel45_Valid_Out & channel25_Kernel45_Valid_Out & channel26_Kernel45_Valid_Out & channel27_Kernel45_Valid_Out & channel28_Kernel45_Valid_Out & channel29_Kernel45_Valid_Out & channel30_Kernel45_Valid_Out & channel31_Kernel45_Valid_Out & channel32_Kernel45_Valid_Out;

	wire channel1_Kernel46_Valid_Out, channel2_Kernel46_Valid_Out, channel3_Kernel46_Valid_Out, channel4_Kernel46_Valid_Out, channel5_Kernel46_Valid_Out, channel6_Kernel46_Valid_Out, channel7_Kernel46_Valid_Out, channel8_Kernel46_Valid_Out, channel9_Kernel46_Valid_Out, channel10_Kernel46_Valid_Out, channel11_Kernel46_Valid_Out, channel12_Kernel46_Valid_Out, channel13_Kernel46_Valid_Out, channel14_Kernel46_Valid_Out, channel15_Kernel46_Valid_Out, channel16_Kernel46_Valid_Out, channel17_Kernel46_Valid_Out, channel18_Kernel46_Valid_Out, channel19_Kernel46_Valid_Out, channel20_Kernel46_Valid_Out, channel21_Kernel46_Valid_Out, channel22_Kernel46_Valid_Out, channel23_Kernel46_Valid_Out, channel24_Kernel46_Valid_Out, channel25_Kernel46_Valid_Out, channel26_Kernel46_Valid_Out, channel27_Kernel46_Valid_Out, channel28_Kernel46_Valid_Out, channel29_Kernel46_Valid_Out, channel30_Kernel46_Valid_Out, channel31_Kernel46_Valid_Out, channel32_Kernel46_Valid_Out;

	assign add_kernel46=channel1_Kernel46_Valid_Out & channel2_Kernel46_Valid_Out & channel3_Kernel46_Valid_Out & channel4_Kernel46_Valid_Out & channel5_Kernel46_Valid_Out & channel6_Kernel46_Valid_Out & channel7_Kernel46_Valid_Out & channel8_Kernel46_Valid_Out & channel9_Kernel46_Valid_Out & channel10_Kernel46_Valid_Out & channel11_Kernel46_Valid_Out & channel12_Kernel46_Valid_Out & channel13_Kernel46_Valid_Out & channel14_Kernel46_Valid_Out & channel15_Kernel46_Valid_Out & channel16_Kernel46_Valid_Out & channel17_Kernel46_Valid_Out & channel18_Kernel46_Valid_Out & channel19_Kernel46_Valid_Out & channel20_Kernel46_Valid_Out & channel21_Kernel46_Valid_Out & channel22_Kernel46_Valid_Out & channel23_Kernel46_Valid_Out & channel24_Kernel46_Valid_Out & channel25_Kernel46_Valid_Out & channel26_Kernel46_Valid_Out & channel27_Kernel46_Valid_Out & channel28_Kernel46_Valid_Out & channel29_Kernel46_Valid_Out & channel30_Kernel46_Valid_Out & channel31_Kernel46_Valid_Out & channel32_Kernel46_Valid_Out;

	wire channel1_Kernel47_Valid_Out, channel2_Kernel47_Valid_Out, channel3_Kernel47_Valid_Out, channel4_Kernel47_Valid_Out, channel5_Kernel47_Valid_Out, channel6_Kernel47_Valid_Out, channel7_Kernel47_Valid_Out, channel8_Kernel47_Valid_Out, channel9_Kernel47_Valid_Out, channel10_Kernel47_Valid_Out, channel11_Kernel47_Valid_Out, channel12_Kernel47_Valid_Out, channel13_Kernel47_Valid_Out, channel14_Kernel47_Valid_Out, channel15_Kernel47_Valid_Out, channel16_Kernel47_Valid_Out, channel17_Kernel47_Valid_Out, channel18_Kernel47_Valid_Out, channel19_Kernel47_Valid_Out, channel20_Kernel47_Valid_Out, channel21_Kernel47_Valid_Out, channel22_Kernel47_Valid_Out, channel23_Kernel47_Valid_Out, channel24_Kernel47_Valid_Out, channel25_Kernel47_Valid_Out, channel26_Kernel47_Valid_Out, channel27_Kernel47_Valid_Out, channel28_Kernel47_Valid_Out, channel29_Kernel47_Valid_Out, channel30_Kernel47_Valid_Out, channel31_Kernel47_Valid_Out, channel32_Kernel47_Valid_Out;

	assign add_kernel47=channel1_Kernel47_Valid_Out & channel2_Kernel47_Valid_Out & channel3_Kernel47_Valid_Out & channel4_Kernel47_Valid_Out & channel5_Kernel47_Valid_Out & channel6_Kernel47_Valid_Out & channel7_Kernel47_Valid_Out & channel8_Kernel47_Valid_Out & channel9_Kernel47_Valid_Out & channel10_Kernel47_Valid_Out & channel11_Kernel47_Valid_Out & channel12_Kernel47_Valid_Out & channel13_Kernel47_Valid_Out & channel14_Kernel47_Valid_Out & channel15_Kernel47_Valid_Out & channel16_Kernel47_Valid_Out & channel17_Kernel47_Valid_Out & channel18_Kernel47_Valid_Out & channel19_Kernel47_Valid_Out & channel20_Kernel47_Valid_Out & channel21_Kernel47_Valid_Out & channel22_Kernel47_Valid_Out & channel23_Kernel47_Valid_Out & channel24_Kernel47_Valid_Out & channel25_Kernel47_Valid_Out & channel26_Kernel47_Valid_Out & channel27_Kernel47_Valid_Out & channel28_Kernel47_Valid_Out & channel29_Kernel47_Valid_Out & channel30_Kernel47_Valid_Out & channel31_Kernel47_Valid_Out & channel32_Kernel47_Valid_Out;

	wire channel1_Kernel48_Valid_Out, channel2_Kernel48_Valid_Out, channel3_Kernel48_Valid_Out, channel4_Kernel48_Valid_Out, channel5_Kernel48_Valid_Out, channel6_Kernel48_Valid_Out, channel7_Kernel48_Valid_Out, channel8_Kernel48_Valid_Out, channel9_Kernel48_Valid_Out, channel10_Kernel48_Valid_Out, channel11_Kernel48_Valid_Out, channel12_Kernel48_Valid_Out, channel13_Kernel48_Valid_Out, channel14_Kernel48_Valid_Out, channel15_Kernel48_Valid_Out, channel16_Kernel48_Valid_Out, channel17_Kernel48_Valid_Out, channel18_Kernel48_Valid_Out, channel19_Kernel48_Valid_Out, channel20_Kernel48_Valid_Out, channel21_Kernel48_Valid_Out, channel22_Kernel48_Valid_Out, channel23_Kernel48_Valid_Out, channel24_Kernel48_Valid_Out, channel25_Kernel48_Valid_Out, channel26_Kernel48_Valid_Out, channel27_Kernel48_Valid_Out, channel28_Kernel48_Valid_Out, channel29_Kernel48_Valid_Out, channel30_Kernel48_Valid_Out, channel31_Kernel48_Valid_Out, channel32_Kernel48_Valid_Out;

	assign add_kernel48=channel1_Kernel48_Valid_Out & channel2_Kernel48_Valid_Out & channel3_Kernel48_Valid_Out & channel4_Kernel48_Valid_Out & channel5_Kernel48_Valid_Out & channel6_Kernel48_Valid_Out & channel7_Kernel48_Valid_Out & channel8_Kernel48_Valid_Out & channel9_Kernel48_Valid_Out & channel10_Kernel48_Valid_Out & channel11_Kernel48_Valid_Out & channel12_Kernel48_Valid_Out & channel13_Kernel48_Valid_Out & channel14_Kernel48_Valid_Out & channel15_Kernel48_Valid_Out & channel16_Kernel48_Valid_Out & channel17_Kernel48_Valid_Out & channel18_Kernel48_Valid_Out & channel19_Kernel48_Valid_Out & channel20_Kernel48_Valid_Out & channel21_Kernel48_Valid_Out & channel22_Kernel48_Valid_Out & channel23_Kernel48_Valid_Out & channel24_Kernel48_Valid_Out & channel25_Kernel48_Valid_Out & channel26_Kernel48_Valid_Out & channel27_Kernel48_Valid_Out & channel28_Kernel48_Valid_Out & channel29_Kernel48_Valid_Out & channel30_Kernel48_Valid_Out & channel31_Kernel48_Valid_Out & channel32_Kernel48_Valid_Out;

	wire channel1_Kernel49_Valid_Out, channel2_Kernel49_Valid_Out, channel3_Kernel49_Valid_Out, channel4_Kernel49_Valid_Out, channel5_Kernel49_Valid_Out, channel6_Kernel49_Valid_Out, channel7_Kernel49_Valid_Out, channel8_Kernel49_Valid_Out, channel9_Kernel49_Valid_Out, channel10_Kernel49_Valid_Out, channel11_Kernel49_Valid_Out, channel12_Kernel49_Valid_Out, channel13_Kernel49_Valid_Out, channel14_Kernel49_Valid_Out, channel15_Kernel49_Valid_Out, channel16_Kernel49_Valid_Out, channel17_Kernel49_Valid_Out, channel18_Kernel49_Valid_Out, channel19_Kernel49_Valid_Out, channel20_Kernel49_Valid_Out, channel21_Kernel49_Valid_Out, channel22_Kernel49_Valid_Out, channel23_Kernel49_Valid_Out, channel24_Kernel49_Valid_Out, channel25_Kernel49_Valid_Out, channel26_Kernel49_Valid_Out, channel27_Kernel49_Valid_Out, channel28_Kernel49_Valid_Out, channel29_Kernel49_Valid_Out, channel30_Kernel49_Valid_Out, channel31_Kernel49_Valid_Out, channel32_Kernel49_Valid_Out;

	assign add_kernel49=channel1_Kernel49_Valid_Out & channel2_Kernel49_Valid_Out & channel3_Kernel49_Valid_Out & channel4_Kernel49_Valid_Out & channel5_Kernel49_Valid_Out & channel6_Kernel49_Valid_Out & channel7_Kernel49_Valid_Out & channel8_Kernel49_Valid_Out & channel9_Kernel49_Valid_Out & channel10_Kernel49_Valid_Out & channel11_Kernel49_Valid_Out & channel12_Kernel49_Valid_Out & channel13_Kernel49_Valid_Out & channel14_Kernel49_Valid_Out & channel15_Kernel49_Valid_Out & channel16_Kernel49_Valid_Out & channel17_Kernel49_Valid_Out & channel18_Kernel49_Valid_Out & channel19_Kernel49_Valid_Out & channel20_Kernel49_Valid_Out & channel21_Kernel49_Valid_Out & channel22_Kernel49_Valid_Out & channel23_Kernel49_Valid_Out & channel24_Kernel49_Valid_Out & channel25_Kernel49_Valid_Out & channel26_Kernel49_Valid_Out & channel27_Kernel49_Valid_Out & channel28_Kernel49_Valid_Out & channel29_Kernel49_Valid_Out & channel30_Kernel49_Valid_Out & channel31_Kernel49_Valid_Out & channel32_Kernel49_Valid_Out;

	wire channel1_Kernel50_Valid_Out, channel2_Kernel50_Valid_Out, channel3_Kernel50_Valid_Out, channel4_Kernel50_Valid_Out, channel5_Kernel50_Valid_Out, channel6_Kernel50_Valid_Out, channel7_Kernel50_Valid_Out, channel8_Kernel50_Valid_Out, channel9_Kernel50_Valid_Out, channel10_Kernel50_Valid_Out, channel11_Kernel50_Valid_Out, channel12_Kernel50_Valid_Out, channel13_Kernel50_Valid_Out, channel14_Kernel50_Valid_Out, channel15_Kernel50_Valid_Out, channel16_Kernel50_Valid_Out, channel17_Kernel50_Valid_Out, channel18_Kernel50_Valid_Out, channel19_Kernel50_Valid_Out, channel20_Kernel50_Valid_Out, channel21_Kernel50_Valid_Out, channel22_Kernel50_Valid_Out, channel23_Kernel50_Valid_Out, channel24_Kernel50_Valid_Out, channel25_Kernel50_Valid_Out, channel26_Kernel50_Valid_Out, channel27_Kernel50_Valid_Out, channel28_Kernel50_Valid_Out, channel29_Kernel50_Valid_Out, channel30_Kernel50_Valid_Out, channel31_Kernel50_Valid_Out, channel32_Kernel50_Valid_Out;

	assign add_kernel50=channel1_Kernel50_Valid_Out & channel2_Kernel50_Valid_Out & channel3_Kernel50_Valid_Out & channel4_Kernel50_Valid_Out & channel5_Kernel50_Valid_Out & channel6_Kernel50_Valid_Out & channel7_Kernel50_Valid_Out & channel8_Kernel50_Valid_Out & channel9_Kernel50_Valid_Out & channel10_Kernel50_Valid_Out & channel11_Kernel50_Valid_Out & channel12_Kernel50_Valid_Out & channel13_Kernel50_Valid_Out & channel14_Kernel50_Valid_Out & channel15_Kernel50_Valid_Out & channel16_Kernel50_Valid_Out & channel17_Kernel50_Valid_Out & channel18_Kernel50_Valid_Out & channel19_Kernel50_Valid_Out & channel20_Kernel50_Valid_Out & channel21_Kernel50_Valid_Out & channel22_Kernel50_Valid_Out & channel23_Kernel50_Valid_Out & channel24_Kernel50_Valid_Out & channel25_Kernel50_Valid_Out & channel26_Kernel50_Valid_Out & channel27_Kernel50_Valid_Out & channel28_Kernel50_Valid_Out & channel29_Kernel50_Valid_Out & channel30_Kernel50_Valid_Out & channel31_Kernel50_Valid_Out & channel32_Kernel50_Valid_Out;

	wire channel1_Kernel51_Valid_Out, channel2_Kernel51_Valid_Out, channel3_Kernel51_Valid_Out, channel4_Kernel51_Valid_Out, channel5_Kernel51_Valid_Out, channel6_Kernel51_Valid_Out, channel7_Kernel51_Valid_Out, channel8_Kernel51_Valid_Out, channel9_Kernel51_Valid_Out, channel10_Kernel51_Valid_Out, channel11_Kernel51_Valid_Out, channel12_Kernel51_Valid_Out, channel13_Kernel51_Valid_Out, channel14_Kernel51_Valid_Out, channel15_Kernel51_Valid_Out, channel16_Kernel51_Valid_Out, channel17_Kernel51_Valid_Out, channel18_Kernel51_Valid_Out, channel19_Kernel51_Valid_Out, channel20_Kernel51_Valid_Out, channel21_Kernel51_Valid_Out, channel22_Kernel51_Valid_Out, channel23_Kernel51_Valid_Out, channel24_Kernel51_Valid_Out, channel25_Kernel51_Valid_Out, channel26_Kernel51_Valid_Out, channel27_Kernel51_Valid_Out, channel28_Kernel51_Valid_Out, channel29_Kernel51_Valid_Out, channel30_Kernel51_Valid_Out, channel31_Kernel51_Valid_Out, channel32_Kernel51_Valid_Out;

	assign add_kernel51=channel1_Kernel51_Valid_Out & channel2_Kernel51_Valid_Out & channel3_Kernel51_Valid_Out & channel4_Kernel51_Valid_Out & channel5_Kernel51_Valid_Out & channel6_Kernel51_Valid_Out & channel7_Kernel51_Valid_Out & channel8_Kernel51_Valid_Out & channel9_Kernel51_Valid_Out & channel10_Kernel51_Valid_Out & channel11_Kernel51_Valid_Out & channel12_Kernel51_Valid_Out & channel13_Kernel51_Valid_Out & channel14_Kernel51_Valid_Out & channel15_Kernel51_Valid_Out & channel16_Kernel51_Valid_Out & channel17_Kernel51_Valid_Out & channel18_Kernel51_Valid_Out & channel19_Kernel51_Valid_Out & channel20_Kernel51_Valid_Out & channel21_Kernel51_Valid_Out & channel22_Kernel51_Valid_Out & channel23_Kernel51_Valid_Out & channel24_Kernel51_Valid_Out & channel25_Kernel51_Valid_Out & channel26_Kernel51_Valid_Out & channel27_Kernel51_Valid_Out & channel28_Kernel51_Valid_Out & channel29_Kernel51_Valid_Out & channel30_Kernel51_Valid_Out & channel31_Kernel51_Valid_Out & channel32_Kernel51_Valid_Out;

	wire channel1_Kernel52_Valid_Out, channel2_Kernel52_Valid_Out, channel3_Kernel52_Valid_Out, channel4_Kernel52_Valid_Out, channel5_Kernel52_Valid_Out, channel6_Kernel52_Valid_Out, channel7_Kernel52_Valid_Out, channel8_Kernel52_Valid_Out, channel9_Kernel52_Valid_Out, channel10_Kernel52_Valid_Out, channel11_Kernel52_Valid_Out, channel12_Kernel52_Valid_Out, channel13_Kernel52_Valid_Out, channel14_Kernel52_Valid_Out, channel15_Kernel52_Valid_Out, channel16_Kernel52_Valid_Out, channel17_Kernel52_Valid_Out, channel18_Kernel52_Valid_Out, channel19_Kernel52_Valid_Out, channel20_Kernel52_Valid_Out, channel21_Kernel52_Valid_Out, channel22_Kernel52_Valid_Out, channel23_Kernel52_Valid_Out, channel24_Kernel52_Valid_Out, channel25_Kernel52_Valid_Out, channel26_Kernel52_Valid_Out, channel27_Kernel52_Valid_Out, channel28_Kernel52_Valid_Out, channel29_Kernel52_Valid_Out, channel30_Kernel52_Valid_Out, channel31_Kernel52_Valid_Out, channel32_Kernel52_Valid_Out;

	assign add_kernel52=channel1_Kernel52_Valid_Out & channel2_Kernel52_Valid_Out & channel3_Kernel52_Valid_Out & channel4_Kernel52_Valid_Out & channel5_Kernel52_Valid_Out & channel6_Kernel52_Valid_Out & channel7_Kernel52_Valid_Out & channel8_Kernel52_Valid_Out & channel9_Kernel52_Valid_Out & channel10_Kernel52_Valid_Out & channel11_Kernel52_Valid_Out & channel12_Kernel52_Valid_Out & channel13_Kernel52_Valid_Out & channel14_Kernel52_Valid_Out & channel15_Kernel52_Valid_Out & channel16_Kernel52_Valid_Out & channel17_Kernel52_Valid_Out & channel18_Kernel52_Valid_Out & channel19_Kernel52_Valid_Out & channel20_Kernel52_Valid_Out & channel21_Kernel52_Valid_Out & channel22_Kernel52_Valid_Out & channel23_Kernel52_Valid_Out & channel24_Kernel52_Valid_Out & channel25_Kernel52_Valid_Out & channel26_Kernel52_Valid_Out & channel27_Kernel52_Valid_Out & channel28_Kernel52_Valid_Out & channel29_Kernel52_Valid_Out & channel30_Kernel52_Valid_Out & channel31_Kernel52_Valid_Out & channel32_Kernel52_Valid_Out;

	wire channel1_Kernel53_Valid_Out, channel2_Kernel53_Valid_Out, channel3_Kernel53_Valid_Out, channel4_Kernel53_Valid_Out, channel5_Kernel53_Valid_Out, channel6_Kernel53_Valid_Out, channel7_Kernel53_Valid_Out, channel8_Kernel53_Valid_Out, channel9_Kernel53_Valid_Out, channel10_Kernel53_Valid_Out, channel11_Kernel53_Valid_Out, channel12_Kernel53_Valid_Out, channel13_Kernel53_Valid_Out, channel14_Kernel53_Valid_Out, channel15_Kernel53_Valid_Out, channel16_Kernel53_Valid_Out, channel17_Kernel53_Valid_Out, channel18_Kernel53_Valid_Out, channel19_Kernel53_Valid_Out, channel20_Kernel53_Valid_Out, channel21_Kernel53_Valid_Out, channel22_Kernel53_Valid_Out, channel23_Kernel53_Valid_Out, channel24_Kernel53_Valid_Out, channel25_Kernel53_Valid_Out, channel26_Kernel53_Valid_Out, channel27_Kernel53_Valid_Out, channel28_Kernel53_Valid_Out, channel29_Kernel53_Valid_Out, channel30_Kernel53_Valid_Out, channel31_Kernel53_Valid_Out, channel32_Kernel53_Valid_Out;

	assign add_kernel53=channel1_Kernel53_Valid_Out & channel2_Kernel53_Valid_Out & channel3_Kernel53_Valid_Out & channel4_Kernel53_Valid_Out & channel5_Kernel53_Valid_Out & channel6_Kernel53_Valid_Out & channel7_Kernel53_Valid_Out & channel8_Kernel53_Valid_Out & channel9_Kernel53_Valid_Out & channel10_Kernel53_Valid_Out & channel11_Kernel53_Valid_Out & channel12_Kernel53_Valid_Out & channel13_Kernel53_Valid_Out & channel14_Kernel53_Valid_Out & channel15_Kernel53_Valid_Out & channel16_Kernel53_Valid_Out & channel17_Kernel53_Valid_Out & channel18_Kernel53_Valid_Out & channel19_Kernel53_Valid_Out & channel20_Kernel53_Valid_Out & channel21_Kernel53_Valid_Out & channel22_Kernel53_Valid_Out & channel23_Kernel53_Valid_Out & channel24_Kernel53_Valid_Out & channel25_Kernel53_Valid_Out & channel26_Kernel53_Valid_Out & channel27_Kernel53_Valid_Out & channel28_Kernel53_Valid_Out & channel29_Kernel53_Valid_Out & channel30_Kernel53_Valid_Out & channel31_Kernel53_Valid_Out & channel32_Kernel53_Valid_Out;

	wire channel1_Kernel54_Valid_Out, channel2_Kernel54_Valid_Out, channel3_Kernel54_Valid_Out, channel4_Kernel54_Valid_Out, channel5_Kernel54_Valid_Out, channel6_Kernel54_Valid_Out, channel7_Kernel54_Valid_Out, channel8_Kernel54_Valid_Out, channel9_Kernel54_Valid_Out, channel10_Kernel54_Valid_Out, channel11_Kernel54_Valid_Out, channel12_Kernel54_Valid_Out, channel13_Kernel54_Valid_Out, channel14_Kernel54_Valid_Out, channel15_Kernel54_Valid_Out, channel16_Kernel54_Valid_Out, channel17_Kernel54_Valid_Out, channel18_Kernel54_Valid_Out, channel19_Kernel54_Valid_Out, channel20_Kernel54_Valid_Out, channel21_Kernel54_Valid_Out, channel22_Kernel54_Valid_Out, channel23_Kernel54_Valid_Out, channel24_Kernel54_Valid_Out, channel25_Kernel54_Valid_Out, channel26_Kernel54_Valid_Out, channel27_Kernel54_Valid_Out, channel28_Kernel54_Valid_Out, channel29_Kernel54_Valid_Out, channel30_Kernel54_Valid_Out, channel31_Kernel54_Valid_Out, channel32_Kernel54_Valid_Out;

	assign add_kernel54=channel1_Kernel54_Valid_Out & channel2_Kernel54_Valid_Out & channel3_Kernel54_Valid_Out & channel4_Kernel54_Valid_Out & channel5_Kernel54_Valid_Out & channel6_Kernel54_Valid_Out & channel7_Kernel54_Valid_Out & channel8_Kernel54_Valid_Out & channel9_Kernel54_Valid_Out & channel10_Kernel54_Valid_Out & channel11_Kernel54_Valid_Out & channel12_Kernel54_Valid_Out & channel13_Kernel54_Valid_Out & channel14_Kernel54_Valid_Out & channel15_Kernel54_Valid_Out & channel16_Kernel54_Valid_Out & channel17_Kernel54_Valid_Out & channel18_Kernel54_Valid_Out & channel19_Kernel54_Valid_Out & channel20_Kernel54_Valid_Out & channel21_Kernel54_Valid_Out & channel22_Kernel54_Valid_Out & channel23_Kernel54_Valid_Out & channel24_Kernel54_Valid_Out & channel25_Kernel54_Valid_Out & channel26_Kernel54_Valid_Out & channel27_Kernel54_Valid_Out & channel28_Kernel54_Valid_Out & channel29_Kernel54_Valid_Out & channel30_Kernel54_Valid_Out & channel31_Kernel54_Valid_Out & channel32_Kernel54_Valid_Out;

	wire channel1_Kernel55_Valid_Out, channel2_Kernel55_Valid_Out, channel3_Kernel55_Valid_Out, channel4_Kernel55_Valid_Out, channel5_Kernel55_Valid_Out, channel6_Kernel55_Valid_Out, channel7_Kernel55_Valid_Out, channel8_Kernel55_Valid_Out, channel9_Kernel55_Valid_Out, channel10_Kernel55_Valid_Out, channel11_Kernel55_Valid_Out, channel12_Kernel55_Valid_Out, channel13_Kernel55_Valid_Out, channel14_Kernel55_Valid_Out, channel15_Kernel55_Valid_Out, channel16_Kernel55_Valid_Out, channel17_Kernel55_Valid_Out, channel18_Kernel55_Valid_Out, channel19_Kernel55_Valid_Out, channel20_Kernel55_Valid_Out, channel21_Kernel55_Valid_Out, channel22_Kernel55_Valid_Out, channel23_Kernel55_Valid_Out, channel24_Kernel55_Valid_Out, channel25_Kernel55_Valid_Out, channel26_Kernel55_Valid_Out, channel27_Kernel55_Valid_Out, channel28_Kernel55_Valid_Out, channel29_Kernel55_Valid_Out, channel30_Kernel55_Valid_Out, channel31_Kernel55_Valid_Out, channel32_Kernel55_Valid_Out;

	assign add_kernel55=channel1_Kernel55_Valid_Out & channel2_Kernel55_Valid_Out & channel3_Kernel55_Valid_Out & channel4_Kernel55_Valid_Out & channel5_Kernel55_Valid_Out & channel6_Kernel55_Valid_Out & channel7_Kernel55_Valid_Out & channel8_Kernel55_Valid_Out & channel9_Kernel55_Valid_Out & channel10_Kernel55_Valid_Out & channel11_Kernel55_Valid_Out & channel12_Kernel55_Valid_Out & channel13_Kernel55_Valid_Out & channel14_Kernel55_Valid_Out & channel15_Kernel55_Valid_Out & channel16_Kernel55_Valid_Out & channel17_Kernel55_Valid_Out & channel18_Kernel55_Valid_Out & channel19_Kernel55_Valid_Out & channel20_Kernel55_Valid_Out & channel21_Kernel55_Valid_Out & channel22_Kernel55_Valid_Out & channel23_Kernel55_Valid_Out & channel24_Kernel55_Valid_Out & channel25_Kernel55_Valid_Out & channel26_Kernel55_Valid_Out & channel27_Kernel55_Valid_Out & channel28_Kernel55_Valid_Out & channel29_Kernel55_Valid_Out & channel30_Kernel55_Valid_Out & channel31_Kernel55_Valid_Out & channel32_Kernel55_Valid_Out;

	wire channel1_Kernel56_Valid_Out, channel2_Kernel56_Valid_Out, channel3_Kernel56_Valid_Out, channel4_Kernel56_Valid_Out, channel5_Kernel56_Valid_Out, channel6_Kernel56_Valid_Out, channel7_Kernel56_Valid_Out, channel8_Kernel56_Valid_Out, channel9_Kernel56_Valid_Out, channel10_Kernel56_Valid_Out, channel11_Kernel56_Valid_Out, channel12_Kernel56_Valid_Out, channel13_Kernel56_Valid_Out, channel14_Kernel56_Valid_Out, channel15_Kernel56_Valid_Out, channel16_Kernel56_Valid_Out, channel17_Kernel56_Valid_Out, channel18_Kernel56_Valid_Out, channel19_Kernel56_Valid_Out, channel20_Kernel56_Valid_Out, channel21_Kernel56_Valid_Out, channel22_Kernel56_Valid_Out, channel23_Kernel56_Valid_Out, channel24_Kernel56_Valid_Out, channel25_Kernel56_Valid_Out, channel26_Kernel56_Valid_Out, channel27_Kernel56_Valid_Out, channel28_Kernel56_Valid_Out, channel29_Kernel56_Valid_Out, channel30_Kernel56_Valid_Out, channel31_Kernel56_Valid_Out, channel32_Kernel56_Valid_Out;

	assign add_kernel56=channel1_Kernel56_Valid_Out & channel2_Kernel56_Valid_Out & channel3_Kernel56_Valid_Out & channel4_Kernel56_Valid_Out & channel5_Kernel56_Valid_Out & channel6_Kernel56_Valid_Out & channel7_Kernel56_Valid_Out & channel8_Kernel56_Valid_Out & channel9_Kernel56_Valid_Out & channel10_Kernel56_Valid_Out & channel11_Kernel56_Valid_Out & channel12_Kernel56_Valid_Out & channel13_Kernel56_Valid_Out & channel14_Kernel56_Valid_Out & channel15_Kernel56_Valid_Out & channel16_Kernel56_Valid_Out & channel17_Kernel56_Valid_Out & channel18_Kernel56_Valid_Out & channel19_Kernel56_Valid_Out & channel20_Kernel56_Valid_Out & channel21_Kernel56_Valid_Out & channel22_Kernel56_Valid_Out & channel23_Kernel56_Valid_Out & channel24_Kernel56_Valid_Out & channel25_Kernel56_Valid_Out & channel26_Kernel56_Valid_Out & channel27_Kernel56_Valid_Out & channel28_Kernel56_Valid_Out & channel29_Kernel56_Valid_Out & channel30_Kernel56_Valid_Out & channel31_Kernel56_Valid_Out & channel32_Kernel56_Valid_Out;

	wire channel1_Kernel57_Valid_Out, channel2_Kernel57_Valid_Out, channel3_Kernel57_Valid_Out, channel4_Kernel57_Valid_Out, channel5_Kernel57_Valid_Out, channel6_Kernel57_Valid_Out, channel7_Kernel57_Valid_Out, channel8_Kernel57_Valid_Out, channel9_Kernel57_Valid_Out, channel10_Kernel57_Valid_Out, channel11_Kernel57_Valid_Out, channel12_Kernel57_Valid_Out, channel13_Kernel57_Valid_Out, channel14_Kernel57_Valid_Out, channel15_Kernel57_Valid_Out, channel16_Kernel57_Valid_Out, channel17_Kernel57_Valid_Out, channel18_Kernel57_Valid_Out, channel19_Kernel57_Valid_Out, channel20_Kernel57_Valid_Out, channel21_Kernel57_Valid_Out, channel22_Kernel57_Valid_Out, channel23_Kernel57_Valid_Out, channel24_Kernel57_Valid_Out, channel25_Kernel57_Valid_Out, channel26_Kernel57_Valid_Out, channel27_Kernel57_Valid_Out, channel28_Kernel57_Valid_Out, channel29_Kernel57_Valid_Out, channel30_Kernel57_Valid_Out, channel31_Kernel57_Valid_Out, channel32_Kernel57_Valid_Out;

	assign add_kernel57=channel1_Kernel57_Valid_Out & channel2_Kernel57_Valid_Out & channel3_Kernel57_Valid_Out & channel4_Kernel57_Valid_Out & channel5_Kernel57_Valid_Out & channel6_Kernel57_Valid_Out & channel7_Kernel57_Valid_Out & channel8_Kernel57_Valid_Out & channel9_Kernel57_Valid_Out & channel10_Kernel57_Valid_Out & channel11_Kernel57_Valid_Out & channel12_Kernel57_Valid_Out & channel13_Kernel57_Valid_Out & channel14_Kernel57_Valid_Out & channel15_Kernel57_Valid_Out & channel16_Kernel57_Valid_Out & channel17_Kernel57_Valid_Out & channel18_Kernel57_Valid_Out & channel19_Kernel57_Valid_Out & channel20_Kernel57_Valid_Out & channel21_Kernel57_Valid_Out & channel22_Kernel57_Valid_Out & channel23_Kernel57_Valid_Out & channel24_Kernel57_Valid_Out & channel25_Kernel57_Valid_Out & channel26_Kernel57_Valid_Out & channel27_Kernel57_Valid_Out & channel28_Kernel57_Valid_Out & channel29_Kernel57_Valid_Out & channel30_Kernel57_Valid_Out & channel31_Kernel57_Valid_Out & channel32_Kernel57_Valid_Out;

	wire channel1_Kernel58_Valid_Out, channel2_Kernel58_Valid_Out, channel3_Kernel58_Valid_Out, channel4_Kernel58_Valid_Out, channel5_Kernel58_Valid_Out, channel6_Kernel58_Valid_Out, channel7_Kernel58_Valid_Out, channel8_Kernel58_Valid_Out, channel9_Kernel58_Valid_Out, channel10_Kernel58_Valid_Out, channel11_Kernel58_Valid_Out, channel12_Kernel58_Valid_Out, channel13_Kernel58_Valid_Out, channel14_Kernel58_Valid_Out, channel15_Kernel58_Valid_Out, channel16_Kernel58_Valid_Out, channel17_Kernel58_Valid_Out, channel18_Kernel58_Valid_Out, channel19_Kernel58_Valid_Out, channel20_Kernel58_Valid_Out, channel21_Kernel58_Valid_Out, channel22_Kernel58_Valid_Out, channel23_Kernel58_Valid_Out, channel24_Kernel58_Valid_Out, channel25_Kernel58_Valid_Out, channel26_Kernel58_Valid_Out, channel27_Kernel58_Valid_Out, channel28_Kernel58_Valid_Out, channel29_Kernel58_Valid_Out, channel30_Kernel58_Valid_Out, channel31_Kernel58_Valid_Out, channel32_Kernel58_Valid_Out;

	assign add_kernel58=channel1_Kernel58_Valid_Out & channel2_Kernel58_Valid_Out & channel3_Kernel58_Valid_Out & channel4_Kernel58_Valid_Out & channel5_Kernel58_Valid_Out & channel6_Kernel58_Valid_Out & channel7_Kernel58_Valid_Out & channel8_Kernel58_Valid_Out & channel9_Kernel58_Valid_Out & channel10_Kernel58_Valid_Out & channel11_Kernel58_Valid_Out & channel12_Kernel58_Valid_Out & channel13_Kernel58_Valid_Out & channel14_Kernel58_Valid_Out & channel15_Kernel58_Valid_Out & channel16_Kernel58_Valid_Out & channel17_Kernel58_Valid_Out & channel18_Kernel58_Valid_Out & channel19_Kernel58_Valid_Out & channel20_Kernel58_Valid_Out & channel21_Kernel58_Valid_Out & channel22_Kernel58_Valid_Out & channel23_Kernel58_Valid_Out & channel24_Kernel58_Valid_Out & channel25_Kernel58_Valid_Out & channel26_Kernel58_Valid_Out & channel27_Kernel58_Valid_Out & channel28_Kernel58_Valid_Out & channel29_Kernel58_Valid_Out & channel30_Kernel58_Valid_Out & channel31_Kernel58_Valid_Out & channel32_Kernel58_Valid_Out;

	wire channel1_Kernel59_Valid_Out, channel2_Kernel59_Valid_Out, channel3_Kernel59_Valid_Out, channel4_Kernel59_Valid_Out, channel5_Kernel59_Valid_Out, channel6_Kernel59_Valid_Out, channel7_Kernel59_Valid_Out, channel8_Kernel59_Valid_Out, channel9_Kernel59_Valid_Out, channel10_Kernel59_Valid_Out, channel11_Kernel59_Valid_Out, channel12_Kernel59_Valid_Out, channel13_Kernel59_Valid_Out, channel14_Kernel59_Valid_Out, channel15_Kernel59_Valid_Out, channel16_Kernel59_Valid_Out, channel17_Kernel59_Valid_Out, channel18_Kernel59_Valid_Out, channel19_Kernel59_Valid_Out, channel20_Kernel59_Valid_Out, channel21_Kernel59_Valid_Out, channel22_Kernel59_Valid_Out, channel23_Kernel59_Valid_Out, channel24_Kernel59_Valid_Out, channel25_Kernel59_Valid_Out, channel26_Kernel59_Valid_Out, channel27_Kernel59_Valid_Out, channel28_Kernel59_Valid_Out, channel29_Kernel59_Valid_Out, channel30_Kernel59_Valid_Out, channel31_Kernel59_Valid_Out, channel32_Kernel59_Valid_Out;

	assign add_kernel59=channel1_Kernel59_Valid_Out & channel2_Kernel59_Valid_Out & channel3_Kernel59_Valid_Out & channel4_Kernel59_Valid_Out & channel5_Kernel59_Valid_Out & channel6_Kernel59_Valid_Out & channel7_Kernel59_Valid_Out & channel8_Kernel59_Valid_Out & channel9_Kernel59_Valid_Out & channel10_Kernel59_Valid_Out & channel11_Kernel59_Valid_Out & channel12_Kernel59_Valid_Out & channel13_Kernel59_Valid_Out & channel14_Kernel59_Valid_Out & channel15_Kernel59_Valid_Out & channel16_Kernel59_Valid_Out & channel17_Kernel59_Valid_Out & channel18_Kernel59_Valid_Out & channel19_Kernel59_Valid_Out & channel20_Kernel59_Valid_Out & channel21_Kernel59_Valid_Out & channel22_Kernel59_Valid_Out & channel23_Kernel59_Valid_Out & channel24_Kernel59_Valid_Out & channel25_Kernel59_Valid_Out & channel26_Kernel59_Valid_Out & channel27_Kernel59_Valid_Out & channel28_Kernel59_Valid_Out & channel29_Kernel59_Valid_Out & channel30_Kernel59_Valid_Out & channel31_Kernel59_Valid_Out & channel32_Kernel59_Valid_Out;

	wire channel1_Kernel60_Valid_Out, channel2_Kernel60_Valid_Out, channel3_Kernel60_Valid_Out, channel4_Kernel60_Valid_Out, channel5_Kernel60_Valid_Out, channel6_Kernel60_Valid_Out, channel7_Kernel60_Valid_Out, channel8_Kernel60_Valid_Out, channel9_Kernel60_Valid_Out, channel10_Kernel60_Valid_Out, channel11_Kernel60_Valid_Out, channel12_Kernel60_Valid_Out, channel13_Kernel60_Valid_Out, channel14_Kernel60_Valid_Out, channel15_Kernel60_Valid_Out, channel16_Kernel60_Valid_Out, channel17_Kernel60_Valid_Out, channel18_Kernel60_Valid_Out, channel19_Kernel60_Valid_Out, channel20_Kernel60_Valid_Out, channel21_Kernel60_Valid_Out, channel22_Kernel60_Valid_Out, channel23_Kernel60_Valid_Out, channel24_Kernel60_Valid_Out, channel25_Kernel60_Valid_Out, channel26_Kernel60_Valid_Out, channel27_Kernel60_Valid_Out, channel28_Kernel60_Valid_Out, channel29_Kernel60_Valid_Out, channel30_Kernel60_Valid_Out, channel31_Kernel60_Valid_Out, channel32_Kernel60_Valid_Out;

	assign add_kernel60=channel1_Kernel60_Valid_Out & channel2_Kernel60_Valid_Out & channel3_Kernel60_Valid_Out & channel4_Kernel60_Valid_Out & channel5_Kernel60_Valid_Out & channel6_Kernel60_Valid_Out & channel7_Kernel60_Valid_Out & channel8_Kernel60_Valid_Out & channel9_Kernel60_Valid_Out & channel10_Kernel60_Valid_Out & channel11_Kernel60_Valid_Out & channel12_Kernel60_Valid_Out & channel13_Kernel60_Valid_Out & channel14_Kernel60_Valid_Out & channel15_Kernel60_Valid_Out & channel16_Kernel60_Valid_Out & channel17_Kernel60_Valid_Out & channel18_Kernel60_Valid_Out & channel19_Kernel60_Valid_Out & channel20_Kernel60_Valid_Out & channel21_Kernel60_Valid_Out & channel22_Kernel60_Valid_Out & channel23_Kernel60_Valid_Out & channel24_Kernel60_Valid_Out & channel25_Kernel60_Valid_Out & channel26_Kernel60_Valid_Out & channel27_Kernel60_Valid_Out & channel28_Kernel60_Valid_Out & channel29_Kernel60_Valid_Out & channel30_Kernel60_Valid_Out & channel31_Kernel60_Valid_Out & channel32_Kernel60_Valid_Out;

	wire channel1_Kernel61_Valid_Out, channel2_Kernel61_Valid_Out, channel3_Kernel61_Valid_Out, channel4_Kernel61_Valid_Out, channel5_Kernel61_Valid_Out, channel6_Kernel61_Valid_Out, channel7_Kernel61_Valid_Out, channel8_Kernel61_Valid_Out, channel9_Kernel61_Valid_Out, channel10_Kernel61_Valid_Out, channel11_Kernel61_Valid_Out, channel12_Kernel61_Valid_Out, channel13_Kernel61_Valid_Out, channel14_Kernel61_Valid_Out, channel15_Kernel61_Valid_Out, channel16_Kernel61_Valid_Out, channel17_Kernel61_Valid_Out, channel18_Kernel61_Valid_Out, channel19_Kernel61_Valid_Out, channel20_Kernel61_Valid_Out, channel21_Kernel61_Valid_Out, channel22_Kernel61_Valid_Out, channel23_Kernel61_Valid_Out, channel24_Kernel61_Valid_Out, channel25_Kernel61_Valid_Out, channel26_Kernel61_Valid_Out, channel27_Kernel61_Valid_Out, channel28_Kernel61_Valid_Out, channel29_Kernel61_Valid_Out, channel30_Kernel61_Valid_Out, channel31_Kernel61_Valid_Out, channel32_Kernel61_Valid_Out;

	assign add_kernel61=channel1_Kernel61_Valid_Out & channel2_Kernel61_Valid_Out & channel3_Kernel61_Valid_Out & channel4_Kernel61_Valid_Out & channel5_Kernel61_Valid_Out & channel6_Kernel61_Valid_Out & channel7_Kernel61_Valid_Out & channel8_Kernel61_Valid_Out & channel9_Kernel61_Valid_Out & channel10_Kernel61_Valid_Out & channel11_Kernel61_Valid_Out & channel12_Kernel61_Valid_Out & channel13_Kernel61_Valid_Out & channel14_Kernel61_Valid_Out & channel15_Kernel61_Valid_Out & channel16_Kernel61_Valid_Out & channel17_Kernel61_Valid_Out & channel18_Kernel61_Valid_Out & channel19_Kernel61_Valid_Out & channel20_Kernel61_Valid_Out & channel21_Kernel61_Valid_Out & channel22_Kernel61_Valid_Out & channel23_Kernel61_Valid_Out & channel24_Kernel61_Valid_Out & channel25_Kernel61_Valid_Out & channel26_Kernel61_Valid_Out & channel27_Kernel61_Valid_Out & channel28_Kernel61_Valid_Out & channel29_Kernel61_Valid_Out & channel30_Kernel61_Valid_Out & channel31_Kernel61_Valid_Out & channel32_Kernel61_Valid_Out;

	wire channel1_Kernel62_Valid_Out, channel2_Kernel62_Valid_Out, channel3_Kernel62_Valid_Out, channel4_Kernel62_Valid_Out, channel5_Kernel62_Valid_Out, channel6_Kernel62_Valid_Out, channel7_Kernel62_Valid_Out, channel8_Kernel62_Valid_Out, channel9_Kernel62_Valid_Out, channel10_Kernel62_Valid_Out, channel11_Kernel62_Valid_Out, channel12_Kernel62_Valid_Out, channel13_Kernel62_Valid_Out, channel14_Kernel62_Valid_Out, channel15_Kernel62_Valid_Out, channel16_Kernel62_Valid_Out, channel17_Kernel62_Valid_Out, channel18_Kernel62_Valid_Out, channel19_Kernel62_Valid_Out, channel20_Kernel62_Valid_Out, channel21_Kernel62_Valid_Out, channel22_Kernel62_Valid_Out, channel23_Kernel62_Valid_Out, channel24_Kernel62_Valid_Out, channel25_Kernel62_Valid_Out, channel26_Kernel62_Valid_Out, channel27_Kernel62_Valid_Out, channel28_Kernel62_Valid_Out, channel29_Kernel62_Valid_Out, channel30_Kernel62_Valid_Out, channel31_Kernel62_Valid_Out, channel32_Kernel62_Valid_Out;

	assign add_kernel62=channel1_Kernel62_Valid_Out & channel2_Kernel62_Valid_Out & channel3_Kernel62_Valid_Out & channel4_Kernel62_Valid_Out & channel5_Kernel62_Valid_Out & channel6_Kernel62_Valid_Out & channel7_Kernel62_Valid_Out & channel8_Kernel62_Valid_Out & channel9_Kernel62_Valid_Out & channel10_Kernel62_Valid_Out & channel11_Kernel62_Valid_Out & channel12_Kernel62_Valid_Out & channel13_Kernel62_Valid_Out & channel14_Kernel62_Valid_Out & channel15_Kernel62_Valid_Out & channel16_Kernel62_Valid_Out & channel17_Kernel62_Valid_Out & channel18_Kernel62_Valid_Out & channel19_Kernel62_Valid_Out & channel20_Kernel62_Valid_Out & channel21_Kernel62_Valid_Out & channel22_Kernel62_Valid_Out & channel23_Kernel62_Valid_Out & channel24_Kernel62_Valid_Out & channel25_Kernel62_Valid_Out & channel26_Kernel62_Valid_Out & channel27_Kernel62_Valid_Out & channel28_Kernel62_Valid_Out & channel29_Kernel62_Valid_Out & channel30_Kernel62_Valid_Out & channel31_Kernel62_Valid_Out & channel32_Kernel62_Valid_Out;

	wire channel1_Kernel63_Valid_Out, channel2_Kernel63_Valid_Out, channel3_Kernel63_Valid_Out, channel4_Kernel63_Valid_Out, channel5_Kernel63_Valid_Out, channel6_Kernel63_Valid_Out, channel7_Kernel63_Valid_Out, channel8_Kernel63_Valid_Out, channel9_Kernel63_Valid_Out, channel10_Kernel63_Valid_Out, channel11_Kernel63_Valid_Out, channel12_Kernel63_Valid_Out, channel13_Kernel63_Valid_Out, channel14_Kernel63_Valid_Out, channel15_Kernel63_Valid_Out, channel16_Kernel63_Valid_Out, channel17_Kernel63_Valid_Out, channel18_Kernel63_Valid_Out, channel19_Kernel63_Valid_Out, channel20_Kernel63_Valid_Out, channel21_Kernel63_Valid_Out, channel22_Kernel63_Valid_Out, channel23_Kernel63_Valid_Out, channel24_Kernel63_Valid_Out, channel25_Kernel63_Valid_Out, channel26_Kernel63_Valid_Out, channel27_Kernel63_Valid_Out, channel28_Kernel63_Valid_Out, channel29_Kernel63_Valid_Out, channel30_Kernel63_Valid_Out, channel31_Kernel63_Valid_Out, channel32_Kernel63_Valid_Out;

	assign add_kernel63=channel1_Kernel63_Valid_Out & channel2_Kernel63_Valid_Out & channel3_Kernel63_Valid_Out & channel4_Kernel63_Valid_Out & channel5_Kernel63_Valid_Out & channel6_Kernel63_Valid_Out & channel7_Kernel63_Valid_Out & channel8_Kernel63_Valid_Out & channel9_Kernel63_Valid_Out & channel10_Kernel63_Valid_Out & channel11_Kernel63_Valid_Out & channel12_Kernel63_Valid_Out & channel13_Kernel63_Valid_Out & channel14_Kernel63_Valid_Out & channel15_Kernel63_Valid_Out & channel16_Kernel63_Valid_Out & channel17_Kernel63_Valid_Out & channel18_Kernel63_Valid_Out & channel19_Kernel63_Valid_Out & channel20_Kernel63_Valid_Out & channel21_Kernel63_Valid_Out & channel22_Kernel63_Valid_Out & channel23_Kernel63_Valid_Out & channel24_Kernel63_Valid_Out & channel25_Kernel63_Valid_Out & channel26_Kernel63_Valid_Out & channel27_Kernel63_Valid_Out & channel28_Kernel63_Valid_Out & channel29_Kernel63_Valid_Out & channel30_Kernel63_Valid_Out & channel31_Kernel63_Valid_Out & channel32_Kernel63_Valid_Out;

	wire channel1_Kernel64_Valid_Out, channel2_Kernel64_Valid_Out, channel3_Kernel64_Valid_Out, channel4_Kernel64_Valid_Out, channel5_Kernel64_Valid_Out, channel6_Kernel64_Valid_Out, channel7_Kernel64_Valid_Out, channel8_Kernel64_Valid_Out, channel9_Kernel64_Valid_Out, channel10_Kernel64_Valid_Out, channel11_Kernel64_Valid_Out, channel12_Kernel64_Valid_Out, channel13_Kernel64_Valid_Out, channel14_Kernel64_Valid_Out, channel15_Kernel64_Valid_Out, channel16_Kernel64_Valid_Out, channel17_Kernel64_Valid_Out, channel18_Kernel64_Valid_Out, channel19_Kernel64_Valid_Out, channel20_Kernel64_Valid_Out, channel21_Kernel64_Valid_Out, channel22_Kernel64_Valid_Out, channel23_Kernel64_Valid_Out, channel24_Kernel64_Valid_Out, channel25_Kernel64_Valid_Out, channel26_Kernel64_Valid_Out, channel27_Kernel64_Valid_Out, channel28_Kernel64_Valid_Out, channel29_Kernel64_Valid_Out, channel30_Kernel64_Valid_Out, channel31_Kernel64_Valid_Out, channel32_Kernel64_Valid_Out;

	assign add_kernel64=channel1_Kernel64_Valid_Out & channel2_Kernel64_Valid_Out & channel3_Kernel64_Valid_Out & channel4_Kernel64_Valid_Out & channel5_Kernel64_Valid_Out & channel6_Kernel64_Valid_Out & channel7_Kernel64_Valid_Out & channel8_Kernel64_Valid_Out & channel9_Kernel64_Valid_Out & channel10_Kernel64_Valid_Out & channel11_Kernel64_Valid_Out & channel12_Kernel64_Valid_Out & channel13_Kernel64_Valid_Out & channel14_Kernel64_Valid_Out & channel15_Kernel64_Valid_Out & channel16_Kernel64_Valid_Out & channel17_Kernel64_Valid_Out & channel18_Kernel64_Valid_Out & channel19_Kernel64_Valid_Out & channel20_Kernel64_Valid_Out & channel21_Kernel64_Valid_Out & channel22_Kernel64_Valid_Out & channel23_Kernel64_Valid_Out & channel24_Kernel64_Valid_Out & channel25_Kernel64_Valid_Out & channel26_Kernel64_Valid_Out & channel27_Kernel64_Valid_Out & channel28_Kernel64_Valid_Out & channel29_Kernel64_Valid_Out & channel30_Kernel64_Valid_Out & channel31_Kernel64_Valid_Out & channel32_Kernel64_Valid_Out;


	wire [31:0] bn1_Data_Out, bn2_Data_Out, bn3_Data_Out, bn4_Data_Out, bn5_Data_Out, bn6_Data_Out, bn7_Data_Out, bn8_Data_Out, bn9_Data_Out, bn10_Data_Out, bn11_Data_Out, bn12_Data_Out, bn13_Data_Out, bn14_Data_Out, bn15_Data_Out, bn16_Data_Out, bn17_Data_Out, bn18_Data_Out, bn19_Data_Out, bn20_Data_Out, bn21_Data_Out, bn22_Data_Out, bn23_Data_Out, bn24_Data_Out, bn25_Data_Out, bn26_Data_Out, bn27_Data_Out, bn28_Data_Out, bn29_Data_Out, bn30_Data_Out, bn31_Data_Out, bn32_Data_Out, bn33_Data_Out, bn34_Data_Out, bn35_Data_Out, bn36_Data_Out, bn37_Data_Out, bn38_Data_Out, bn39_Data_Out, bn40_Data_Out, bn41_Data_Out, bn42_Data_Out, bn43_Data_Out, bn44_Data_Out, bn45_Data_Out, bn46_Data_Out, bn47_Data_Out, bn48_Data_Out, bn49_Data_Out, bn50_Data_Out, bn51_Data_Out, bn52_Data_Out, bn53_Data_Out, bn54_Data_Out, bn55_Data_Out, bn56_Data_Out, bn57_Data_Out, bn58_Data_Out, bn59_Data_Out, bn60_Data_Out, bn61_Data_Out, bn62_Data_Out, bn63_Data_Out, bn64_Data_Out;

	wire bn1_Valid_Out, bn2_Valid_Out, bn3_Valid_Out, bn4_Valid_Out, bn5_Valid_Out, bn6_Valid_Out, bn7_Valid_Out, bn8_Valid_Out, bn9_Valid_Out, bn10_Valid_Out, bn11_Valid_Out, bn12_Valid_Out, bn13_Valid_Out, bn14_Valid_Out, bn15_Valid_Out, bn16_Valid_Out, bn17_Valid_Out, bn18_Valid_Out, bn19_Valid_Out, bn20_Valid_Out, bn21_Valid_Out, bn22_Valid_Out, bn23_Valid_Out, bn24_Valid_Out, bn25_Valid_Out, bn26_Valid_Out, bn27_Valid_Out, bn28_Valid_Out, bn29_Valid_Out, bn30_Valid_Out, bn31_Valid_Out, bn32_Valid_Out, bn33_Valid_Out, bn34_Valid_Out, bn35_Valid_Out, bn36_Valid_Out, bn37_Valid_Out, bn38_Valid_Out, bn39_Valid_Out, bn40_Valid_Out, bn41_Valid_Out, bn42_Valid_Out, bn43_Valid_Out, bn44_Valid_Out, bn45_Valid_Out, bn46_Valid_Out, bn47_Valid_Out, bn48_Valid_Out, bn49_Valid_Out, bn50_Valid_Out, bn51_Valid_Out, bn52_Valid_Out, bn53_Valid_Out, bn54_Valid_Out, bn55_Valid_Out, bn56_Valid_Out, bn57_Valid_Out, bn58_Valid_Out, bn59_Valid_Out, bn60_Valid_Out, bn61_Valid_Out, bn62_Valid_Out, bn63_Valid_Out, bn64_Valid_Out;

	wire rl1_Valid_Out, rl2_Valid_Out, rl3_Valid_Out, rl4_Valid_Out, rl5_Valid_Out, rl6_Valid_Out, rl7_Valid_Out, rl8_Valid_Out, rl9_Valid_Out, rl10_Valid_Out, rl11_Valid_Out, rl12_Valid_Out, rl13_Valid_Out, rl14_Valid_Out, rl15_Valid_Out, rl16_Valid_Out, rl17_Valid_Out, rl18_Valid_Out, rl19_Valid_Out, rl20_Valid_Out, rl21_Valid_Out, rl22_Valid_Out, rl23_Valid_Out, rl24_Valid_Out, rl25_Valid_Out, rl26_Valid_Out, rl27_Valid_Out, rl28_Valid_Out, rl29_Valid_Out, rl30_Valid_Out, rl31_Valid_Out, rl32_Valid_Out, rl33_Valid_Out, rl34_Valid_Out, rl35_Valid_Out, rl36_Valid_Out, rl37_Valid_Out, rl38_Valid_Out, rl39_Valid_Out, rl40_Valid_Out, rl41_Valid_Out, rl42_Valid_Out, rl43_Valid_Out, rl44_Valid_Out, rl45_Valid_Out, rl46_Valid_Out, rl47_Valid_Out, rl48_Valid_Out, rl49_Valid_Out, rl50_Valid_Out, rl51_Valid_Out, rl52_Valid_Out, rl53_Valid_Out, rl54_Valid_Out, rl55_Valid_Out, rl56_Valid_Out, rl57_Valid_Out, rl58_Valid_Out, rl59_Valid_Out, rl60_Valid_Out, rl61_Valid_Out, rl62_Valid_Out, rl63_Valid_Out, rl64_Valid_Out;

	 assign Valid_Out = rl1_Valid_Out & rl2_Valid_Out & rl3_Valid_Out & rl4_Valid_Out & rl5_Valid_Out & rl6_Valid_Out & rl7_Valid_Out & rl8_Valid_Out & rl9_Valid_Out & rl10_Valid_Out & rl11_Valid_Out & rl12_Valid_Out & rl13_Valid_Out & rl14_Valid_Out & rl15_Valid_Out & rl16_Valid_Out & rl17_Valid_Out & rl18_Valid_Out & rl19_Valid_Out & rl20_Valid_Out & rl21_Valid_Out & rl22_Valid_Out & rl23_Valid_Out & rl24_Valid_Out & rl25_Valid_Out & rl26_Valid_Out & rl27_Valid_Out & rl28_Valid_Out & rl29_Valid_Out & rl30_Valid_Out & rl31_Valid_Out & rl32_Valid_Out & rl33_Valid_Out & rl34_Valid_Out & rl35_Valid_Out & rl36_Valid_Out & rl37_Valid_Out & rl38_Valid_Out & rl39_Valid_Out & rl40_Valid_Out & rl41_Valid_Out & rl42_Valid_Out & rl43_Valid_Out & rl44_Valid_Out & rl45_Valid_Out & rl46_Valid_Out & rl47_Valid_Out & rl48_Valid_Out & rl49_Valid_Out & rl50_Valid_Out & rl51_Valid_Out & rl52_Valid_Out & rl53_Valid_Out & rl54_Valid_Out & rl55_Valid_Out & rl56_Valid_Out & rl57_Valid_Out & rl58_Valid_Out & rl59_Valid_Out & rl60_Valid_Out & rl61_Valid_Out & rl62_Valid_Out & rl63_Valid_Out & rl64_Valid_Out;
//////////KERNEL1//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111110110001010011010011101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110100111000011010011000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110110100111011100101010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111101010001011101000010010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111110111101010001010001000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110000100000111001011100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111111000010011111101000101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111110000011111110101011001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111110111110001111000000100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110001001010111001011000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111111011110001010000101011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111110101001111111000111011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111101111111110011011001101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111101111001100010100011001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111101001101110101100001001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111110101100010100110000010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111110110111011111111000101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111110010110111111001010000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111110100111001000001100100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110011011011011000010011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111111001110101101101001010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111100000100011100010000010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111100101000100011011010011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111111000100111111011100000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111110001010100011000011010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111110101100101100000000101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111111000000010000010010111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111111000011111011110010001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111110000001111001110101111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110101111110111010010001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111101110110111100000010111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel1_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel1 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110110001100110100100101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel1[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel1_Valid_Out)
	);
	Adder_32input add_k1(
		.Data1(Data_Out_Kernel1[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel1[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel1[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel1[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel1[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel1[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel1[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel1[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel1[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel1[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel1[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel1[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel1[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel1[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel1[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel1[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel1[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel1[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel1[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel1[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel1[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel1[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel1[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel1[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel1[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel1[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel1[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel1[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel1[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel1[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel1[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel1[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel1),
		.Data_Out(add_k1_Data_Out),
		.Valid_Out(add_kernel1_Valid_Out)
	);
	Batch_Norm bn_kernel1(
		.Data_A(32'b00111110100011110111100111101010),
		.Data_B(32'b10111110101111010101011111001001),
		.Data_In(add_k1_Data_Out),
		.Valid_In(add_kernel1_Valid_Out),
		.Data_Out(bn1_Data_Out),
		.Valid_Out(bn1_Valid_Out)
	);
	Relu_Core rl_kernel1(
		.Data_In(bn1_Data_Out),
		.Valid_In(bn1_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT-1:0]),
		.Valid_Out(rl1_Valid_Out)
	);
//////////KERNEL2//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111101110011000011111000111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111101110011111100000101100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111101110010111010011011011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111100110010000111000110101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111110110010010110111111010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111110101110000100100111100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111110111011001000001000100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111110100000001011100000110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111011101001010111000100001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111111000010011101001110011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111101001111010111000001100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111111001000000011100111111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111101111101001001111000101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111111000100010000010101010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111111010011000111000110010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111111001100100011100000001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111110100100000100110110111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111111000010000010010100110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110100000001100101111110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111110101001100001111011010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111111000110011110101001111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111110010111101001110000001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110111100001011110110010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111101101001100001000100011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111110000010000000000011111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110000011001001111101000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110101101001100100001011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110110111111001101111110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111110001010011100001011010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110011011100010111010011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111110101101000110100001100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel2_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel2 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110011011100001101001011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel2[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel2_Valid_Out)
	);
	Adder_32input add_k2(
		.Data1(Data_Out_Kernel2[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel2[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel2[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel2[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel2[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel2[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel2[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel2[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel2[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel2[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel2[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel2[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel2[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel2[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel2[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel2[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel2[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel2[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel2[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel2[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel2[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel2[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel2[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel2[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel2[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel2[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel2[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel2[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel2[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel2[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel2[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel2[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel2),
		.Data_Out(add_k2_Data_Out),
		.Valid_Out(add_kernel2_Valid_Out)
	);
	Batch_Norm bn_kernel2(
		.Data_A(32'b00111110010011101100101111111100),
		.Data_B(32'b10111101111001101011101110100010),
		.Data_In(add_k2_Data_Out),
		.Valid_In(add_kernel2_Valid_Out),
		.Data_Out(bn2_Data_Out),
		.Valid_Out(bn2_Valid_Out)
	);
	Relu_Core rl_kernel2(
		.Data_In(bn2_Data_Out),
		.Valid_In(bn2_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Valid_Out(rl2_Valid_Out)
	);
//////////KERNEL3//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111101010011011000010011000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111110101110101101110000100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110011001010110001010100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110100011110000001111111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111110111001101100000001101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111101010101001000110100111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111110000010111011001110001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111110101111001100001010001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111111001100101101000010101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111110011001101110101011100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111110010111001101111011101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110010001000100110011101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111101100000110011001000110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111110000001000100100001101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111100011010011010001111000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111111010100110011010011010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111100110001010110100011101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111110111111011110110010010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111111010010101110110000010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111110111110100110101010011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111100010010001111011101111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111111000101110000110110011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111101011100100001110010001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111100011101000111001000110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111111000000100111010001101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111111001101100111110010100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110000111110110001110100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111101101010101011101110111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111110011110111100000000101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111111000101010100010110000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111110100001111000011110111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel3_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel3 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111110010000011001000001111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel3[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel3_Valid_Out)
	);
	Adder_32input add_k3(
		.Data1(Data_Out_Kernel3[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel3[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel3[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel3[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel3[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel3[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel3[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel3[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel3[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel3[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel3[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel3[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel3[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel3[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel3[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel3[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel3[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel3[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel3[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel3[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel3[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel3[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel3[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel3[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel3[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel3[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel3[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel3[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel3[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel3[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel3[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel3[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel3),
		.Data_Out(add_k3_Data_Out),
		.Valid_Out(add_kernel3_Valid_Out)
	);
	Batch_Norm bn_kernel3(
		.Data_A(32'b00111110100000000010100101100110),
		.Data_B(32'b00111101010011101000101111101010),
		.Data_In(add_k3_Data_Out),
		.Valid_In(add_kernel3_Valid_Out),
		.Data_Out(bn3_Data_Out),
		.Valid_Out(bn3_Valid_Out)
	);
	Relu_Core rl_kernel3(
		.Data_In(bn3_Data_Out),
		.Valid_In(bn3_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(rl3_Valid_Out)
	);
//////////KERNEL4//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111110110100011100110111110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111110001101000011100101001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110000110001101110100011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111111000110101111101100011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111110110001110010101010000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111110110011100010000000010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111110010111110101110011110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111110110100111101100100111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111111010001000110001111010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110101001111010010000101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111110010110110010111100100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111101111110110111010010001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111101111110011000000001000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111110001101111001010011010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110111100111010010001010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111110110110011001101101010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111101100010001010101011011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111111000101010010110100110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111110000101011110000100110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111110101110000010110101010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111111001000001001110000100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111111000100001010001010111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111111001000111001011001000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111101111010100111011011101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111110011011101010110011110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111101101101101101100111010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111101101110010111110101101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111101000000001111111100111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111101110011001000111101010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110011000111001101011100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111110100100010000111100111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel4_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel4 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111110100101001110111110001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel4[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel4_Valid_Out)
	);
	Adder_32input add_k4(
		.Data1(Data_Out_Kernel4[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel4[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel4[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel4[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel4[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel4[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel4[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel4[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel4[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel4[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel4[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel4[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel4[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel4[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel4[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel4[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel4[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel4[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel4[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel4[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel4[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel4[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel4[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel4[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel4[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel4[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel4[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel4[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel4[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel4[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel4[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel4[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel4),
		.Data_Out(add_k4_Data_Out),
		.Valid_Out(add_kernel4_Valid_Out)
	);
	Batch_Norm bn_kernel4(
		.Data_A(32'b00111110011110111110010011000001),
		.Data_B(32'b10111111000011100101101001000010),
		.Data_In(add_k4_Data_Out),
		.Valid_In(add_kernel4_Valid_Out),
		.Data_Out(bn4_Data_Out),
		.Valid_Out(bn4_Valid_Out)
	);
	Relu_Core rl_kernel4(
		.Data_In(bn4_Data_Out),
		.Valid_In(bn4_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(rl4_Valid_Out)
	);
//////////KERNEL5//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111001110011100000010100100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111101101010010001001111101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110001110110101110001011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110101011010110000100010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111110000011101010001101011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110111101100111001000110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111111000010011111010100110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111101000100010000010001111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111110001111101000101000101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111111001110101110101010001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110100110101000000111011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111110101001011011011011000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111110111111101011111110111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111110100001010101111101111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111101111101101100101100010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111101110110100001011111101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111110101001101001110000100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111111000010011010110111001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111101100000010111100000110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111110111111011111000101100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110001010111010110001101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111111001000011111110110011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111100100111110110100111000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111101000110110010000010100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111111001111010100101011110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111110101001010010010111100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111111000100011001110110100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111100010001100101010101011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111110111110101010110111101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111101000111010001100001000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111101011110111001010010010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel5_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel5 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111110011100001110001001111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel5[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel5_Valid_Out)
	);
	Adder_32input add_k5(
		.Data1(Data_Out_Kernel5[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel5[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel5[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel5[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel5[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel5[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel5[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel5[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel5[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel5[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel5[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel5[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel5[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel5[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel5[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel5[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel5[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel5[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel5[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel5[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel5[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel5[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel5[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel5[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel5[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel5[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel5[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel5[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel5[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel5[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel5[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel5[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel5),
		.Data_Out(add_k5_Data_Out),
		.Valid_Out(add_kernel5_Valid_Out)
	);
	Batch_Norm bn_kernel5(
		.Data_A(32'b00111110100001001110100110001011),
		.Data_B(32'b00111111000011000110011011111111),
		.Data_In(add_k5_Data_Out),
		.Valid_In(add_kernel5_Valid_Out),
		.Data_Out(bn5_Data_Out),
		.Valid_Out(bn5_Valid_Out)
	);
	Relu_Core rl_kernel5(
		.Data_In(bn5_Data_Out),
		.Valid_In(bn5_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(rl5_Valid_Out)
	);
//////////KERNEL6//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110101010011111011010011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111010110101010101011110011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111111000101101101100001011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110001110111111101110011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111101100100001110111100111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111111000101011011001010111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111110011011011000101101110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111111000010010101100110001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111101110001101011011010001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111110100110100110101001101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110100001000101110010001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110000100000101110000011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111100110001010011011100100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111110011011110110001000011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111101010110100011010111111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111111001011011101111111101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110000111110110100110011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110111011000010110000111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111110111011011111010010100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111100111101011100010001011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110110100110110010010011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111110101110011010010111111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110100000001010111101110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111101011100001101001001101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111111100010101100101110100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110001111000001100101000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111110100011001110101000110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111110001011011000111001101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111110001011011100101110011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111101110101011011000000010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111110010100101110010101010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel6_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel6 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110111101101011011110110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel6[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel6_Valid_Out)
	);
	Adder_32input add_k6(
		.Data1(Data_Out_Kernel6[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel6[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel6[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel6[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel6[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel6[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel6[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel6[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel6[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel6[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel6[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel6[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel6[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel6[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel6[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel6[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel6[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel6[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel6[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel6[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel6[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel6[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel6[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel6[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel6[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel6[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel6[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel6[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel6[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel6[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel6[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel6[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel6),
		.Data_Out(add_k6_Data_Out),
		.Valid_Out(add_kernel6_Valid_Out)
	);
	Batch_Norm bn_kernel6(
		.Data_A(32'b00111110011011010001101111101011),
		.Data_B(32'b00111110011000110010110000101011),
		.Data_In(add_k6_Data_Out),
		.Valid_In(add_kernel6_Valid_Out),
		.Data_Out(bn6_Data_Out),
		.Valid_Out(bn6_Valid_Out)
	);
	Relu_Core rl_kernel6(
		.Data_In(bn6_Data_Out),
		.Valid_In(bn6_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(rl6_Valid_Out)
	);
//////////KERNEL7//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110100000000000111001000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111111000101000001110001000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110001110101101001011101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110100111001001100100101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111110100000011001000010111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111110110110110110110010010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111110001101110111111111111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111110110111110101111011011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110000000100111010111111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111111001010100110010101001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110110111111010011001011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111101100111110011101010001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111101110100001101111011011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111011110000111111000111111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110100100100010101100110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111111000100001110101100001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111110100000100100001010110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111111000101000110000011110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110111101111000100010010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111110001001000011101001000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110100011110110011100110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111110111001110010011101001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110000001001001010101011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111101111110011011011000000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111110001110111000001110010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110100101001010011010001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111111000011111001000000100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111111010000011000001010000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111110000001010010000000010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111110011100111111010110101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111111001111011100110111010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel7_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel7 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111110100000011000111101100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel7[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel7_Valid_Out)
	);
	Adder_32input add_k7(
		.Data1(Data_Out_Kernel7[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel7[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel7[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel7[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel7[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel7[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel7[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel7[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel7[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel7[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel7[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel7[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel7[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel7[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel7[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel7[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel7[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel7[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel7[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel7[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel7[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel7[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel7[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel7[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel7[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel7[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel7[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel7[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel7[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel7[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel7[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel7[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel7),
		.Data_Out(add_k7_Data_Out),
		.Valid_Out(add_kernel7_Valid_Out)
	);
	Batch_Norm bn_kernel7(
		.Data_A(32'b00111110100000011101000101100111),
		.Data_B(32'b10111101100101111111111111000000),
		.Data_In(add_k7_Data_Out),
		.Valid_In(add_kernel7_Valid_Out),
		.Data_Out(bn7_Data_Out),
		.Valid_Out(bn7_Valid_Out)
	);
	Relu_Core rl_kernel7(
		.Data_In(bn7_Data_Out),
		.Valid_In(bn7_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(rl7_Valid_Out)
	);
//////////KERNEL8//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111101011110011001010111101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111110101001010100011101110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110101101011011011111000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111101100000001010101111111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111110101011100101010111110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110001010111100111110011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111101101001110010101110011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111110101111101010010011010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110101001001110000100100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111111001001000111010011100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111101011001010011110010110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110100000100011110101101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111101111011110100000010100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111111000010110101111000010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110111101001010001111111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111110101000100111010111110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110001110011100100101100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110101100100111011111100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111111001000100010011111010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111110101011011101111000100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111101110010011101001111111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111110001100011101000101001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111111001001101100010110000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111101100001011110111010011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111110100110111101000110000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111110100011101111101100101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111110101010101100001111110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111111101011001000101010000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111101110110101011100010110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110101101000010011111011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111101110111101001110001110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel8_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel8 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111101010010110000110000001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel8[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel8_Valid_Out)
	);
	Adder_32input add_k8(
		.Data1(Data_Out_Kernel8[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel8[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel8[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel8[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel8[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel8[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel8[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel8[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel8[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel8[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel8[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel8[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel8[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel8[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel8[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel8[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel8[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel8[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel8[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel8[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel8[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel8[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel8[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel8[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel8[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel8[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel8[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel8[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel8[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel8[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel8[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel8[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel8),
		.Data_Out(add_k8_Data_Out),
		.Valid_Out(add_kernel8_Valid_Out)
	);
	Batch_Norm bn_kernel8(
		.Data_A(32'b00111110100100011111011010101111),
		.Data_B(32'b00111110100110010101101111111010),
		.Data_In(add_k8_Data_Out),
		.Valid_In(add_kernel8_Valid_Out),
		.Data_Out(bn8_Data_Out),
		.Valid_Out(bn8_Valid_Out)
	);
	Relu_Core rl_kernel8(
		.Data_In(bn8_Data_Out),
		.Valid_In(bn8_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(rl8_Valid_Out)
	);
//////////KERNEL9//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111100100110110011001110100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111101101110000110010010111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110101011101101101101110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110110110011000111110110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111110111011100000110100101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110001001010011011110001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111110001101110100101011011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111110001010110101000110100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110111100011111011111110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110101011101000010010000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111111000000100100111111110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110100010100010000100010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111111100001010011011101110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111101001110100111110110111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110010110010001111001101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111110110001011110100111001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111101111001111000011110110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111110110110011001000101110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111101100011110011001111011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110000001000001100101010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110100001001111010010001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111110110101110101110100101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111110110111010011101000000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111101100101101111111010011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111111100000001100110101010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111110101101001101101001111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111110000110110001011110011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110110001111110100100011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111110010100101000010000101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111101111110111111111000001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111110001001100110110011001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel9_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel9 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110111000011011110000010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel9[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel9_Valid_Out)
	);
	Adder_32input add_k9(
		.Data1(Data_Out_Kernel9[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel9[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel9[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel9[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel9[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel9[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel9[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel9[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel9[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel9[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel9[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel9[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel9[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel9[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel9[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel9[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel9[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel9[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel9[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel9[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel9[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel9[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel9[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel9[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel9[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel9[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel9[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel9[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel9[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel9[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel9[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel9[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel9),
		.Data_Out(add_k9_Data_Out),
		.Valid_Out(add_kernel9_Valid_Out)
	);
	Batch_Norm bn_kernel9(
		.Data_A(32'b00111110010101110000000101101001),
		.Data_B(32'b00111110100110011000101100100011),
		.Data_In(add_k9_Data_Out),
		.Valid_In(add_kernel9_Valid_Out),
		.Data_Out(bn9_Data_Out),
		.Valid_Out(bn9_Valid_Out)
	);
	Relu_Core rl_kernel9(
		.Data_In(bn9_Data_Out),
		.Valid_In(bn9_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(rl9_Valid_Out)
	);
//////////KERNEL10//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111100001011111010111101110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110000110001000011111000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111111001000001010110001110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110001110001010100100100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111110110010010111011001011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111101001010101001111111110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111111001001110111011111001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111110100110011111100111101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111111001010100100100011100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111101011111111001011100110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111101011110101100100101100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111101100001111101110000000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111100000010100110000100101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111101110100110101100101111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111111001110001000000111001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111100010001110100100000001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111111000000101010010101001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111111011011111101001001100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110100100000011010110001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111111001100110001010110010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111111001000111000100101100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111101110010001001011111111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110100000010001000010100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111100110010011111010000001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111110000001111011010001001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111011010010001000000110111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111101001001001011010011101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111111000000001010001100101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111110010001110001101011011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111111000110111111001000100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111101000111001111001100111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel10_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel10 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111110000011001010111100010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel10[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel10_Valid_Out)
	);
	Adder_32input add_k10(
		.Data1(Data_Out_Kernel10[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel10[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel10[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel10[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel10[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel10[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel10[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel10[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel10[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel10[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel10[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel10[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel10[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel10[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel10[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel10[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel10[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel10[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel10[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel10[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel10[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel10[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel10[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel10[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel10[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel10[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel10[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel10[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel10[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel10[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel10[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel10[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel10),
		.Data_Out(add_k10_Data_Out),
		.Valid_Out(add_kernel10_Valid_Out)
	);
	Batch_Norm bn_kernel10(
		.Data_A(32'b00111110011011000000110110101110),
		.Data_B(32'b00111111000101000110010101100010),
		.Data_In(add_k10_Data_Out),
		.Valid_In(add_kernel10_Valid_Out),
		.Data_Out(bn10_Data_Out),
		.Valid_Out(bn10_Valid_Out)
	);
	Relu_Core rl_kernel10(
		.Data_In(bn10_Data_Out),
		.Valid_In(bn10_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(rl10_Valid_Out)
	);
//////////KERNEL11//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111110111010100101010001000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111101110100110100011111011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110010100000100100111101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111101111101011100000000111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111110010101110011000001110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111110111010011000101110101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111111001011101100001001100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111110101000111011110100111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111110001111011101111111001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111111010010100001100000000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111110101110001100011110000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111101100010001000101000111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111111010010001101111100011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111110000100010011000000100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110100010110011110011011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111110010101101001110001101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111110000000111011010000110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111110100110110010011101110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110001100100111011100011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110111011101111000100000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110100001110011000111001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111110010011101001011010010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111110110010011100010000110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111111001010110011101101110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111110100001001110101011101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111101001000110111010000100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111111000000011111111010010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110100111000100011000110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111101110110100100001000011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111110110101000010110011001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111111011001100011101000100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel11_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel11 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111101001101011010100110010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel11[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel11_Valid_Out)
	);
	Adder_32input add_k11(
		.Data1(Data_Out_Kernel11[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel11[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel11[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel11[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel11[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel11[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel11[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel11[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel11[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel11[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel11[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel11[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel11[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel11[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel11[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel11[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel11[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel11[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel11[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel11[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel11[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel11[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel11[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel11[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel11[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel11[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel11[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel11[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel11[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel11[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel11[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel11[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel11),
		.Data_Out(add_k11_Data_Out),
		.Valid_Out(add_kernel11_Valid_Out)
	);
	Batch_Norm bn_kernel11(
		.Data_A(32'b00111110011011110011011111111111),
		.Data_B(32'b10111101001001111111101001011001),
		.Data_In(add_k11_Data_Out),
		.Valid_In(add_kernel11_Valid_Out),
		.Data_Out(bn11_Data_Out),
		.Valid_Out(bn11_Valid_Out)
	);
	Relu_Core rl_kernel11(
		.Data_In(bn11_Data_Out),
		.Valid_In(bn11_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(rl11_Valid_Out)
	);
//////////KERNEL12//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111110001000110000101110000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111111010111110010011011000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110110011000100000000101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111101000010000110100010011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111110011100101010101000010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111101110010101111011111110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111110100111101000001101111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111110010000111001010101001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111110010001001101111011001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110110000101100001111101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110010110101100110111001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111111000110101000000000100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111111000001100100100000111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111110110010001100101110111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110011011011011110000101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111110010101111000010011110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111100001100111000011000010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111100001110110001001011110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110000101010111110000010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111110100001010110111010001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111100110110010111110000010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111110011010101101111011001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110001000001100000000110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111111000100001101011010101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111110101001010100111111100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110110110100111011110000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111111000000100110001110111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111110100011011010111001111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111111000111110111011101100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111110000100001010110000011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111111000000011100101001001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel12_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel12 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111110101100010010000000110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel12[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel12_Valid_Out)
	);
	Adder_32input add_k12(
		.Data1(Data_Out_Kernel12[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel12[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel12[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel12[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel12[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel12[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel12[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel12[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel12[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel12[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel12[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel12[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel12[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel12[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel12[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel12[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel12[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel12[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel12[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel12[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel12[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel12[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel12[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel12[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel12[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel12[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel12[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel12[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel12[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel12[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel12[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel12[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel12),
		.Data_Out(add_k12_Data_Out),
		.Valid_Out(add_kernel12_Valid_Out)
	);
	Batch_Norm bn_kernel12(
		.Data_A(32'b00111110011000101000101111111001),
		.Data_B(32'b00111110010011100110110010111000),
		.Data_In(add_k12_Data_Out),
		.Valid_In(add_kernel12_Valid_Out),
		.Data_Out(bn12_Data_Out),
		.Valid_Out(bn12_Valid_Out)
	);
	Relu_Core rl_kernel12(
		.Data_In(bn12_Data_Out),
		.Valid_In(bn12_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(rl12_Valid_Out)
	);
//////////KERNEL13//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111110110010000111100101010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111101010101101011010001011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111111000110001001011000010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110110011110010010000001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111110000101111000011000000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111101111010101100001010001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111110010001001111000101010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111011100101000010000100000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111100010110101110001011011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111101111110110010010101111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111110100110001110111100001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111111000011010111101110010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111101111111110010000010111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111111011101101011101001001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110101111010100011010000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111110110010000000111000110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111111000000010000010110101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111110101010100110110001001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110001100000110011111110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111110000010110000010111101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111100111101011101101100000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111110100101001001000101101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111101101100011110111011001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111110100101001100101011010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111110110001101111111000001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111101011110101000100001000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111111000000110011001001100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111101000011000100011110101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111111001001100110011010100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111101010101100101011100011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111101111001111101110110010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel13_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel13 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110110111100000111011111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel13[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel13_Valid_Out)
	);
	Adder_32input add_k13(
		.Data1(Data_Out_Kernel13[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel13[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel13[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel13[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel13[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel13[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel13[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel13[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel13[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel13[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel13[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel13[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel13[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel13[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel13[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel13[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel13[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel13[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel13[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel13[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel13[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel13[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel13[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel13[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel13[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel13[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel13[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel13[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel13[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel13[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel13[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel13[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel13),
		.Data_Out(add_k13_Data_Out),
		.Valid_Out(add_kernel13_Valid_Out)
	);
	Batch_Norm bn_kernel13(
		.Data_A(32'b00111110100000110011011000000110),
		.Data_B(32'b10111111100110001111111011000000),
		.Data_In(add_k13_Data_Out),
		.Valid_In(add_kernel13_Valid_Out),
		.Data_Out(bn13_Data_Out),
		.Valid_Out(bn13_Valid_Out)
	);
	Relu_Core rl_kernel13(
		.Data_In(bn13_Data_Out),
		.Valid_In(bn13_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(rl13_Valid_Out)
	);
//////////KERNEL14//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111110111001001010001001001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110101100110011101001100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110101100111111011001110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111111000000111001100100000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111101110010111100011001010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110100100101101011100011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111101001101010101110110101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111101101000110010111111101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110111000110000011100100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111111001001111001111001001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111110001101111111110101101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110001000011110001111111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111111001111101011110101001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111110000111010000100010101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110111100100001010010010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111101001010011001100111110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110000110001111111111010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111110110110101011000111000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111111000101111010000110001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110100010000000011101001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111111010000101000101101110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111110110010100000100100100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111110010111101101001011001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111110100010001010011110010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111110001100001110111011001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111110100011111110001100011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111110111011000010101110010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111101101101000110011011100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111110110001100111110101010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111110101111110011100101010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111101000000100101000111111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel14_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel14 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111110110001010010101110000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel14[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel14_Valid_Out)
	);
	Adder_32input add_k14(
		.Data1(Data_Out_Kernel14[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel14[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel14[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel14[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel14[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel14[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel14[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel14[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel14[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel14[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel14[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel14[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel14[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel14[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel14[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel14[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel14[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel14[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel14[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel14[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel14[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel14[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel14[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel14[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel14[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel14[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel14[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel14[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel14[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel14[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel14[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel14[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel14),
		.Data_Out(add_k14_Data_Out),
		.Valid_Out(add_kernel14_Valid_Out)
	);
	Batch_Norm bn_kernel14(
		.Data_A(32'b00111110011111110000011010010100),
		.Data_B(32'b00111110110100000100000001111110),
		.Data_In(add_k14_Data_Out),
		.Valid_In(add_kernel14_Valid_Out),
		.Data_Out(bn14_Data_Out),
		.Valid_Out(bn14_Valid_Out)
	);
	Relu_Core rl_kernel14(
		.Data_In(bn14_Data_Out),
		.Valid_In(bn14_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(rl14_Valid_Out)
	);
//////////KERNEL15//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110100101101010001110111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111111000110000100000000001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111111000010001010011110011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110010001110101110011000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111101100100000100111100110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111110100000101011011111110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111110110111101001000000101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111111000000101000000010110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110110000000101110110000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111110101010110001001000010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111111001101001101111010111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110100111111001101001111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111110001111101101000111001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111110100111110100110000001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110011111100101011100000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111101011100100000010010110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111110011111101100001010000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111100111101000101011111110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110011011011111110000111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111111000011100010011101000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111111000100000001000100000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111110110000000100011000000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111110010011110011000010110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111111010100000010011010111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111110001100100100011011101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111110010011110100010110111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111110100100011101101101111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110011001110000000111011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111110000100111101110101110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111111000100001111100001111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111110100000101111111010000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel15_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel15 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110101110110101001111000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel15[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel15_Valid_Out)
	);
	Adder_32input add_k15(
		.Data1(Data_Out_Kernel15[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel15[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel15[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel15[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel15[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel15[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel15[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel15[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel15[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel15[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel15[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel15[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel15[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel15[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel15[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel15[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel15[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel15[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel15[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel15[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel15[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel15[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel15[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel15[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel15[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel15[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel15[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel15[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel15[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel15[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel15[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel15[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel15),
		.Data_Out(add_k15_Data_Out),
		.Valid_Out(add_kernel15_Valid_Out)
	);
	Batch_Norm bn_kernel15(
		.Data_A(32'b00111110100010001100110010101101),
		.Data_B(32'b00111110101110010101110100001110),
		.Data_In(add_k15_Data_Out),
		.Valid_In(add_kernel15_Valid_Out),
		.Data_Out(bn15_Data_Out),
		.Valid_Out(bn15_Valid_Out)
	);
	Relu_Core rl_kernel15(
		.Data_In(bn15_Data_Out),
		.Valid_In(bn15_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(rl15_Valid_Out)
	);
//////////KERNEL16//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110110000001101000101101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111111000101010110010110111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111101100000011101111000100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110100100001000101011010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111111001010101101011001010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111110000011001101011111001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111101000001010000011110101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111110100100010110000011100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111101100111001100001100101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111110011001010100001001010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110111001111011001010001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111111001100100111000101111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111101111010001101000011011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111110100001101101111001100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110100110000001000001111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111110101110011000001001100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110110100101111001000001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110011011000110011000100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111110100101111011101110001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110010111111100010100110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110101110011110111010100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111110000011000010010011110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111110001001001001000100011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111110110010110000000111110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111110011001101100101001001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111110110001100000111000011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111110101001111011001110101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110010110000111101100011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111111010010011100110011110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110010100101111011010110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111101111000010000110100110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel16_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel16 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111110100000001111100000101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel16[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel16_Valid_Out)
	);
	Adder_32input add_k16(
		.Data1(Data_Out_Kernel16[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel16[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel16[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel16[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel16[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel16[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel16[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel16[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel16[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel16[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel16[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel16[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel16[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel16[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel16[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel16[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel16[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel16[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel16[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel16[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel16[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel16[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel16[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel16[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel16[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel16[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel16[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel16[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel16[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel16[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel16[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel16[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel16),
		.Data_Out(add_k16_Data_Out),
		.Valid_Out(add_kernel16_Valid_Out)
	);
	Batch_Norm bn_kernel16(
		.Data_A(32'b00111110010110110101110010100111),
		.Data_B(32'b00111111001011001001000011101000),
		.Data_In(add_k16_Data_Out),
		.Valid_In(add_kernel16_Valid_Out),
		.Data_Out(bn16_Data_Out),
		.Valid_Out(bn16_Valid_Out)
	);
	Relu_Core rl_kernel16(
		.Data_In(bn16_Data_Out),
		.Valid_In(bn16_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(rl16_Valid_Out)
	);
//////////KERNEL17//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110111001001111000101101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110110010110011000011110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111101110000111100011111000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111101111001100010011010110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111110101011010001001111001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111111000100001101000011100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111111000100110011111110011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111110100101110101110011100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111110100110110010000111011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110101101111110110010111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110100111100111111001000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110011111110001110100000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110110000101001110001000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111110111111010001100011110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110100110000110111111001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111100101111111000101111011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110000100101110101111011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111110101100111001101110100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111111000101111001010000010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111101101001101011111011010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111111000111101101111010100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111110001000001001011101101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111110011100010000001100001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111110100101100101000011001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111111000110100011101001110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110111100100100100100001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110101111101010011100001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111110010001101101010011101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111110000110110100010000011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111111001001101100011111100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111110101001010101100100101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel17_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel17 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111110011111001001111101111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel17[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel17_Valid_Out)
	);
	Adder_32input add_k17(
		.Data1(Data_Out_Kernel17[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel17[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel17[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel17[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel17[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel17[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel17[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel17[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel17[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel17[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel17[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel17[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel17[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel17[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel17[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel17[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel17[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel17[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel17[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel17[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel17[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel17[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel17[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel17[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel17[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel17[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel17[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel17[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel17[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel17[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel17[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel17[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel17),
		.Data_Out(add_k17_Data_Out),
		.Valid_Out(add_kernel17_Valid_Out)
	);
	Batch_Norm bn_kernel17(
		.Data_A(32'b00111110011000001010010101110001),
		.Data_B(32'b00111110111111010111101000100101),
		.Data_In(add_k17_Data_Out),
		.Valid_In(add_kernel17_Valid_Out),
		.Data_Out(bn17_Data_Out),
		.Valid_Out(bn17_Valid_Out)
	);
	Relu_Core rl_kernel17(
		.Data_In(bn17_Data_Out),
		.Valid_In(bn17_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(rl17_Valid_Out)
	);
//////////KERNEL18//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111101010011011100111011111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111111011100001001111111101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111111000110010110001010110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111101101100101010001100001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111101111100101111010110111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111110110011010110111001100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111111010010010011010101101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111101110000001101100010100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111110111101101010110101000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111010101111100110001001110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111101110100110010101110001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111110101011010000101111100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111100011111010100110010100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111101001110001000000101001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111101001001001011111110011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111111000011100101001110011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110101011001011111001001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111101101100011101000111011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110000101111110011010001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111111001010010000100100101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110100011000100011100100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111110101010101100101110011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111101001001110111111000110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111110111010110111011011111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111101011011000000001011010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111111001000000001100100010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111110101101111101001110001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111101100001001011111100100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111110010110001110111001010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111110111110101001011001001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111101110000100110101000010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel18_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel18 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111101100000011101111001001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel18[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel18_Valid_Out)
	);
	Adder_32input add_k18(
		.Data1(Data_Out_Kernel18[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel18[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel18[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel18[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel18[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel18[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel18[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel18[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel18[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel18[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel18[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel18[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel18[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel18[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel18[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel18[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel18[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel18[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel18[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel18[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel18[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel18[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel18[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel18[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel18[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel18[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel18[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel18[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel18[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel18[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel18[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel18[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel18),
		.Data_Out(add_k18_Data_Out),
		.Valid_Out(add_kernel18_Valid_Out)
	);
	Batch_Norm bn_kernel18(
		.Data_A(32'b00111110100000101111011101011010),
		.Data_B(32'b10111110010110110100010001000111),
		.Data_In(add_k18_Data_Out),
		.Valid_In(add_kernel18_Valid_Out),
		.Data_Out(bn18_Data_Out),
		.Valid_Out(bn18_Valid_Out)
	);
	Relu_Core rl_kernel18(
		.Data_In(bn18_Data_Out),
		.Valid_In(bn18_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(rl18_Valid_Out)
	);
//////////KERNEL19//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111110100110101101001100001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111101111001100100110000000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111101001010011011101110000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110110100011101100010100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111111010110110011101011001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110001010010010101011101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111110010010110100101100101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111101111010000000011100011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111101010010011010111001110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111110000001101111101100010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111110010100111100010101001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110001110000010111011100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110010011001001100001010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111011111100111011010001000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111111000110010010000000101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111111001100000100000000110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110101010110101001111111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111110111001000111100100101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111101011010011001000010010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111101011101001001110011111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111101011101001000111110011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111011111010101101000100111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111110010101100110110001110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111111000000110011010111101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111101011110011111101110100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111111000010011101110111000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110001100111110111101101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110010010111011000111010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111111001001111010101000001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111111000000001101101011000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111110101011010100100100011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel19_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel19 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111110110011111101111001001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel19[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel19_Valid_Out)
	);
	Adder_32input add_k19(
		.Data1(Data_Out_Kernel19[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel19[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel19[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel19[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel19[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel19[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel19[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel19[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel19[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel19[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel19[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel19[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel19[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel19[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel19[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel19[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel19[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel19[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel19[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel19[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel19[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel19[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel19[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel19[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel19[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel19[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel19[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel19[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel19[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel19[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel19[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel19[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel19),
		.Data_Out(add_k19_Data_Out),
		.Valid_Out(add_kernel19_Valid_Out)
	);
	Batch_Norm bn_kernel19(
		.Data_A(32'b00111110100010000011000010110100),
		.Data_B(32'b10111111100001001101000000100111),
		.Data_In(add_k19_Data_Out),
		.Valid_In(add_kernel19_Valid_Out),
		.Data_Out(bn19_Data_Out),
		.Valid_Out(bn19_Valid_Out)
	);
	Relu_Core rl_kernel19(
		.Data_In(bn19_Data_Out),
		.Valid_In(bn19_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(rl19_Valid_Out)
	);
//////////KERNEL20//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111110111111001010101100010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111101101111111110011110011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110111000011000000010011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111100110000011100011110110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111101001010110110111011011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111101111010100110111000100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111101110001110011000110010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111110110111110101011101010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110011101111101010010011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111110001000111100101100111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111101000000110111011011111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111111001100100010101101100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110010000001101011111101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111111011111010011111101011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110000100101011010101111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111110100101011001110111111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110011110001011000111010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111110100000101101000110000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111101000111011111001101010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110100111011101100011000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110000010111000100100101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111101010011010100101011110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111110000111001101101100110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111110100001111111110010011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111110000011011110101111100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111111001100101001111011000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110011110110011100101111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111101001011011011011001101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111110100101000010001111101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111111010011111101101100111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111111000000101100010010000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel20_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel20 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110000101101010110010001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel20[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel20_Valid_Out)
	);
	Adder_32input add_k20(
		.Data1(Data_Out_Kernel20[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel20[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel20[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel20[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel20[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel20[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel20[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel20[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel20[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel20[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel20[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel20[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel20[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel20[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel20[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel20[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel20[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel20[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel20[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel20[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel20[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel20[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel20[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel20[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel20[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel20[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel20[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel20[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel20[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel20[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel20[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel20[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel20),
		.Data_Out(add_k20_Data_Out),
		.Valid_Out(add_kernel20_Valid_Out)
	);
	Batch_Norm bn_kernel20(
		.Data_A(32'b00111110011100001010011011010010),
		.Data_B(32'b10111111001111011111011100110001),
		.Data_In(add_k20_Data_Out),
		.Valid_In(add_kernel20_Valid_Out),
		.Data_Out(bn20_Data_Out),
		.Valid_Out(bn20_Valid_Out)
	);
	Relu_Core rl_kernel20(
		.Data_In(bn20_Data_Out),
		.Valid_In(bn20_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(rl20_Valid_Out)
	);
//////////KERNEL21//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110101001010001011011101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110111010000001001010001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110100010111000111100111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111111001011100110110100110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111101111001110001000001011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111101001110100010011010101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111110100101000001110010101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111110100100000010111011011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111110101001000100111110001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110010110000000011101111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110100010110101000000011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111111001111110101101001000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111111000000110001101110011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111110101110100100010111011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111101011101000101101110010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111110010001110010000101101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111101110101011000001110101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110100100110001010010111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110101000101001111101110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111111000111001100010000001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111101010111001011001101101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111110100010101001010010101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110101111001000001100000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111110001010010111110010010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111111001110110000100010100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111111000100100101010001101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111101011010101001001110001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111101011100010101100001111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111110011000101001010101000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111110111010100101111000111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111110011110100001001111111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel21_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel21 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111111000001011101100010011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel21[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel21_Valid_Out)
	);
	Adder_32input add_k21(
		.Data1(Data_Out_Kernel21[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel21[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel21[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel21[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel21[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel21[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel21[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel21[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel21[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel21[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel21[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel21[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel21[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel21[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel21[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel21[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel21[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel21[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel21[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel21[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel21[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel21[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel21[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel21[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel21[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel21[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel21[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel21[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel21[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel21[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel21[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel21[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel21),
		.Data_Out(add_k21_Data_Out),
		.Valid_Out(add_kernel21_Valid_Out)
	);
	Batch_Norm bn_kernel21(
		.Data_A(32'b00111110010110101010011011001000),
		.Data_B(32'b00111111010001010111011001001011),
		.Data_In(add_k21_Data_Out),
		.Valid_In(add_kernel21_Valid_Out),
		.Data_Out(bn21_Data_Out),
		.Valid_Out(bn21_Valid_Out)
	);
	Relu_Core rl_kernel21(
		.Data_In(bn21_Data_Out),
		.Valid_In(bn21_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(rl21_Valid_Out)
	);
//////////KERNEL22//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110111101111100011010100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111101111101110011110001111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111111000101001111011100101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110001001001100000101001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111111000111110010110000011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110110110010110000100010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111111000111001011100000000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111110101110000101111100000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110110100001100110110010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111101000011001111001001010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111111001101101010001110110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111111000001001100011101000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111110000101101011010101111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111110101110110110100011001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110010011001111110100011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111110010001000101000000111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110100011011001110011101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110000000001110100011000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110010101010001011101101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111110100000000000100001101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111111000000001011010011111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111110010111001011000010001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111110100001101011100010001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111111000011001111111110101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111111001011101111001011100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111110010011110110011000101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111110100011111110000110110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111101001110011100011010110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111110001000110101001110010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111110000111000001011010010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111101101101000101000000001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel22_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel22 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111110111101011001010000011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel22[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel22_Valid_Out)
	);
	Adder_32input add_k22(
		.Data1(Data_Out_Kernel22[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel22[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel22[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel22[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel22[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel22[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel22[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel22[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel22[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel22[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel22[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel22[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel22[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel22[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel22[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel22[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel22[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel22[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel22[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel22[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel22[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel22[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel22[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel22[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel22[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel22[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel22[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel22[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel22[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel22[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel22[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel22[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel22),
		.Data_Out(add_k22_Data_Out),
		.Valid_Out(add_kernel22_Valid_Out)
	);
	Batch_Norm bn_kernel22(
		.Data_A(32'b00111110011110100100001110000001),
		.Data_B(32'b10111110101010011110110001110000),
		.Data_In(add_k22_Data_Out),
		.Valid_In(add_kernel22_Valid_Out),
		.Data_Out(bn22_Data_Out),
		.Valid_Out(bn22_Valid_Out)
	);
	Relu_Core rl_kernel22(
		.Data_In(bn22_Data_Out),
		.Valid_In(bn22_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(rl22_Valid_Out)
	);
//////////KERNEL23//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111110001110100000000010001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111101100100110111111000110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110100010010101010001011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111101000110010101100000111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111111000000100000011000001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111111001010010101010100111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111101111111011111001000111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111111000001111011101010010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111101111011010110000011010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110010010000100100011111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110100001111110100000000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111110100011001011111111111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111111000101100001110011111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111110100101011101001111001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111100111001010110010011011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111111000001101000011000001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111110101010100110111101100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111111010000100100111000110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111110011000110110101100111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111101101110010011111110010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110010010111011110110110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111110010001000111011100111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111101110001101101000011110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111101000110101001110000111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111110100110011011000010000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111011011010101110001000110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111111000100111011111111010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111111001010000111011101011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111111000000001100101110110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110000110010101101101001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111110000011100010010101100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel23_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel23 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111111000110101111011010100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel23[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel23_Valid_Out)
	);
	Adder_32input add_k23(
		.Data1(Data_Out_Kernel23[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel23[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel23[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel23[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel23[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel23[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel23[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel23[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel23[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel23[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel23[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel23[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel23[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel23[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel23[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel23[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel23[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel23[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel23[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel23[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel23[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel23[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel23[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel23[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel23[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel23[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel23[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel23[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel23[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel23[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel23[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel23[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel23),
		.Data_Out(add_k23_Data_Out),
		.Valid_Out(add_kernel23_Valid_Out)
	);
	Batch_Norm bn_kernel23(
		.Data_A(32'b00111110100001100100000111110010),
		.Data_B(32'b10111110110001100110101110100110),
		.Data_In(add_k23_Data_Out),
		.Valid_In(add_kernel23_Valid_Out),
		.Data_Out(bn23_Data_Out),
		.Valid_Out(bn23_Valid_Out)
	);
	Relu_Core rl_kernel23(
		.Data_In(bn23_Data_Out),
		.Valid_In(bn23_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(rl23_Valid_Out)
	);
//////////KERNEL24//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111101001111011100111100000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111110010111001100011001000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110000100111000011000110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110111101100001101010000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111101110101111011001110110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111110100111011000001011101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111101000111010111010011101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111110110000011110100010111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110010110011000111011010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110101001001111111101110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111111011100100101110010010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111111000000110100111010111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111101011101110111100111111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111110010111011010110111010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110101010111100000101000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111101001010011000010000110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110110010101001010010010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111110001000011110110101001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110111101111001101010011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111110101100101010101110010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110111001101111110110111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111110001011110100000110100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111111010000110000001100100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111111000010111011110011001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111110110010100000110001100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111100100101011100100011000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110101000010011001101100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111101001011000001110011111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111110100001000011000111000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111110111100101011100011101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111110010010011011000000001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel24_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel24 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111110110101010110010001110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel24[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel24_Valid_Out)
	);
	Adder_32input add_k24(
		.Data1(Data_Out_Kernel24[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel24[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel24[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel24[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel24[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel24[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel24[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel24[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel24[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel24[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel24[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel24[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel24[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel24[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel24[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel24[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel24[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel24[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel24[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel24[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel24[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel24[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel24[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel24[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel24[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel24[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel24[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel24[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel24[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel24[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel24[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel24[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel24),
		.Data_Out(add_k24_Data_Out),
		.Valid_Out(add_kernel24_Valid_Out)
	);
	Batch_Norm bn_kernel24(
		.Data_A(32'b00111110011011111100010111101110),
		.Data_B(32'b00111111101000011111110001101110),
		.Data_In(add_k24_Data_Out),
		.Valid_In(add_kernel24_Valid_Out),
		.Data_Out(bn24_Data_Out),
		.Valid_Out(bn24_Valid_Out)
	);
	Relu_Core rl_kernel24(
		.Data_In(bn24_Data_Out),
		.Valid_In(bn24_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(rl24_Valid_Out)
	);
//////////KERNEL25//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111110010110111011101010001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110100101001000111011011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111101100111000111101011100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111101010111000000100101110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111110011000100001001101000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111101001100000110001011010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111111011000011000001001110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111111000100101101101011001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111111001111010101000011010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111110101101110011011101101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111111000011000010001010011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111110110000011001110011000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111110001001000100010010110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111101010110111111011010011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111101110111001100111011100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111101010011101100000000000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111100101111001011101100011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110110111011011101010001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111101101011101110000001000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111100001011101001010110100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110011000100011010101100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111110100110101100111111011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111111000110100101110101110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111110111111111100100100000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111110100100100101101101001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110010110011001000110111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111110011000010100011000010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110110110111001101110010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111101001011101001110000000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111111000001001011011110000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111101010110001010000101011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel25_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel25 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111111001101101111011011111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel25[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel25_Valid_Out)
	);
	Adder_32input add_k25(
		.Data1(Data_Out_Kernel25[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel25[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel25[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel25[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel25[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel25[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel25[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel25[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel25[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel25[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel25[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel25[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel25[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel25[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel25[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel25[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel25[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel25[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel25[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel25[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel25[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel25[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel25[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel25[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel25[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel25[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel25[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel25[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel25[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel25[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel25[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel25[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel25),
		.Data_Out(add_k25_Data_Out),
		.Valid_Out(add_kernel25_Valid_Out)
	);
	Batch_Norm bn_kernel25(
		.Data_A(32'b00111110100001001101101111010101),
		.Data_B(32'b00111110100000101011000100011110),
		.Data_In(add_k25_Data_Out),
		.Valid_In(add_kernel25_Valid_Out),
		.Data_Out(bn25_Data_Out),
		.Valid_Out(bn25_Valid_Out)
	);
	Relu_Core rl_kernel25(
		.Data_In(bn25_Data_Out),
		.Valid_In(bn25_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(rl25_Valid_Out)
	);
//////////KERNEL26//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110110101001100101001000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111111001110011001000010011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110110101001011010001101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111111000111100110011010001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111101111011001101101111011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110110101111011100101100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111110010101101000100100100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111110110011101001101100100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111111000001010000011101100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111111000100000101001101011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110000101010110110110010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111101101110000010110101000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111111001000101011100100110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111100001010010000101000100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110101011100001101101010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111110000111000110010011101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111110011110100011011011100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110100100010110110100100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111101100100111011111010011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111100100000011000001010000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111010100000011011100100001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111111000111101111011111101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111111000000100000101000000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111101101010000011001001010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111110101101101011001001001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111101111010011000101010111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111110000100001111100101100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110000011101010110100111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111101100110111000001110010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110100011100001110001110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111101101100000101110001000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel26_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel26 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111111000000100001001001000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel26[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel26_Valid_Out)
	);
	Adder_32input add_k26(
		.Data1(Data_Out_Kernel26[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel26[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel26[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel26[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel26[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel26[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel26[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel26[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel26[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel26[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel26[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel26[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel26[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel26[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel26[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel26[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel26[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel26[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel26[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel26[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel26[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel26[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel26[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel26[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel26[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel26[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel26[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel26[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel26[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel26[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel26[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel26[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel26),
		.Data_Out(add_k26_Data_Out),
		.Valid_Out(add_kernel26_Valid_Out)
	);
	Batch_Norm bn_kernel26(
		.Data_A(32'b00111110011110111001101010001111),
		.Data_B(32'b00111111011100000000101001101010),
		.Data_In(add_k26_Data_Out),
		.Valid_In(add_kernel26_Valid_Out),
		.Data_Out(bn26_Data_Out),
		.Valid_Out(bn26_Valid_Out)
	);
	Relu_Core rl_kernel26(
		.Data_In(bn26_Data_Out),
		.Valid_In(bn26_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(rl26_Valid_Out)
	);
//////////KERNEL27//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111110110100110001000010010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110110101011000110010010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111101100111011110000010010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111111000000111001010010011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111110000001100100001101101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111110010111110001000100101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111101110001110111010010001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111111001100111110000111111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111110000111111111101110000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111111000101100110000010001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110100100010100000101010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111101110010110101010110111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111111001110000011111101001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111110000000000001101100001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111101001110110001011011010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111111011000110111000101101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110110000100000001101000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110101100010010100011111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110111111000001100010001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110110111111110100000100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110111000111011011000010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111110100010000111100101110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111110010100010010000010111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111100110111011011111010001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111111000101101100001100110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111110010001010000110101111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111110011101100010110011000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111110010110000011000001000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111110111100000100100000011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111100000001101001000110110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111110000101001000110101010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel27_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel27 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111101011000011111110011000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel27[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel27_Valid_Out)
	);
	Adder_32input add_k27(
		.Data1(Data_Out_Kernel27[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel27[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel27[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel27[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel27[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel27[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel27[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel27[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel27[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel27[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel27[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel27[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel27[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel27[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel27[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel27[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel27[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel27[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel27[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel27[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel27[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel27[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel27[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel27[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel27[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel27[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel27[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel27[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel27[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel27[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel27[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel27[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel27),
		.Data_Out(add_k27_Data_Out),
		.Valid_Out(add_kernel27_Valid_Out)
	);
	Batch_Norm bn_kernel27(
		.Data_A(32'b00111110010110101011101001101100),
		.Data_B(32'b10111111000001001011010111101111),
		.Data_In(add_k27_Data_Out),
		.Valid_In(add_kernel27_Valid_Out),
		.Data_Out(bn27_Data_Out),
		.Valid_Out(bn27_Valid_Out)
	);
	Relu_Core rl_kernel27(
		.Data_In(bn27_Data_Out),
		.Valid_In(bn27_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(rl27_Valid_Out)
	);
//////////KERNEL28//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111110000000010010111011111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111110100010010000100010000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110000110000110110010110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110111011101100100011000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111110101101001100101101001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111110000011001111000111100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111110011101111000110111001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111101001101010101011010111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111101000000001011010010011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110100011100000011010101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111101010011001110110100011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111111100000010101111111001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111110110101111000111010100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111110001011001000111001101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110111100100101110101111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111111000101101111010101010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111110111101101110111110101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111101001110100101110011111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110101111101001000001111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110000111111100111010101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110111011000101011000010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111111000010010111110011110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111111001110110101011101001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111110011110110010011011001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111011100001010001011000110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111110110001010110001111101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111101100011010100011001100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111110110111001010010000100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111110100011110010111101000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111100001010011001111111101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111110011100101001110111101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel28_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel28 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110100100101011000111101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel28[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel28_Valid_Out)
	);
	Adder_32input add_k28(
		.Data1(Data_Out_Kernel28[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel28[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel28[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel28[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel28[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel28[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel28[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel28[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel28[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel28[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel28[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel28[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel28[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel28[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel28[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel28[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel28[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel28[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel28[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel28[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel28[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel28[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel28[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel28[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel28[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel28[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel28[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel28[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel28[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel28[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel28[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel28[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel28),
		.Data_Out(add_k28_Data_Out),
		.Valid_Out(add_kernel28_Valid_Out)
	);
	Batch_Norm bn_kernel28(
		.Data_A(32'b00111110100000100011011111101001),
		.Data_B(32'b10111110110100110100111101111010),
		.Data_In(add_k28_Data_Out),
		.Valid_In(add_kernel28_Valid_Out),
		.Data_Out(bn28_Data_Out),
		.Valid_Out(bn28_Valid_Out)
	);
	Relu_Core rl_kernel28(
		.Data_In(bn28_Data_Out),
		.Valid_In(bn28_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(rl28_Valid_Out)
	);
//////////KERNEL29//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111101000010011001100111111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111111100011011011101100010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111101110101010011111110111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111101011100110111011110110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111101101010011111100101111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111110101010111100000001100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111111000001011110110101010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111111000100010111111100000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111101011000000110001000110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110110111111100011111000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110000000111010111011010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111111000100001000010010111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110010010110010001010110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111111000001001100000001100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111111000110000100100010110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111110101110000010011001001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111101100001111000010101111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110101101101100001001110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111101100000111000100111001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111111000001001111110110101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110101001110011101010110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111110100010000001000101101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111101111010010100100110101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111110001101001001001111000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111110011110001111010101000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111110011011111111100001001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111110101101111100011100100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111101101001110111110111101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111110101010011101000001011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111100100000111100100011100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111110101100000101000001011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel29_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel29 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111110011111000100001111100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel29[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel29_Valid_Out)
	);
	Adder_32input add_k29(
		.Data1(Data_Out_Kernel29[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel29[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel29[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel29[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel29[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel29[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel29[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel29[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel29[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel29[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel29[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel29[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel29[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel29[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel29[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel29[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel29[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel29[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel29[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel29[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel29[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel29[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel29[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel29[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel29[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel29[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel29[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel29[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel29[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel29[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel29[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel29[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel29),
		.Data_Out(add_k29_Data_Out),
		.Valid_Out(add_kernel29_Valid_Out)
	);
	Batch_Norm bn_kernel29(
		.Data_A(32'b00111110011111111110000100010101),
		.Data_B(32'b00111111001101010101110011011000),
		.Data_In(add_k29_Data_Out),
		.Valid_In(add_kernel29_Valid_Out),
		.Data_Out(bn29_Data_Out),
		.Valid_Out(bn29_Valid_Out)
	);
	Relu_Core rl_kernel29(
		.Data_In(bn29_Data_Out),
		.Valid_In(bn29_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(rl29_Valid_Out)
	);
//////////KERNEL30//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111101110000010010001101000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110010011000000010010100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110111000011100111110100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111111001111011111110011100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111111001100110111100101101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111111001101000011100011011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111101111011001111100011000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111011101111000100010011111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110111010100000100100011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111110101001110111001001000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111110011101111001010000010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111101111100111001111111110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111101111101111001000000001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111100111101100100011100110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110101010000000000110101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111101101010001010110111110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110111100011010001000111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110110010000001110110001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110111100011111100100111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110001110101000001011111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110100000110110101110011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111100001110111111010001001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110001010100001111110001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111101011111011001100001000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111111000010000110001000011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111110110001110100001011011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110100000101011011100101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111111000011100011101110110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111101100000100011110111001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111101011110101100111000100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111110101110000000000001000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel30_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel30 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111010000011110010011001011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel30[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel30_Valid_Out)
	);
	Adder_32input add_k30(
		.Data1(Data_Out_Kernel30[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel30[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel30[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel30[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel30[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel30[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel30[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel30[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel30[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel30[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel30[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel30[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel30[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel30[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel30[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel30[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel30[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel30[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel30[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel30[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel30[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel30[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel30[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel30[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel30[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel30[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel30[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel30[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel30[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel30[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel30[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel30[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel30),
		.Data_Out(add_k30_Data_Out),
		.Valid_Out(add_kernel30_Valid_Out)
	);
	Batch_Norm bn_kernel30(
		.Data_A(32'b00111110011111100100111010000011),
		.Data_B(32'b10111111100000111011000000011101),
		.Data_In(add_k30_Data_Out),
		.Valid_In(add_kernel30_Valid_Out),
		.Data_Out(bn30_Data_Out),
		.Valid_Out(bn30_Valid_Out)
	);
	Relu_Core rl_kernel30(
		.Data_In(bn30_Data_Out),
		.Valid_In(bn30_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(rl30_Valid_Out)
	);
//////////KERNEL31//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111110100010011111011011111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111011110001101101000000101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110010001001000100110010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111111000010110111111001001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111110111110011110111011010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111100111011000001001111101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111101110101001100111110101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111100110110000001111100001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111110111100110101010011001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111110101001011100001011011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111110101111000101001101101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111111000011100100111100001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111101100010101100110100011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111110000100100101010001101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111111000010101101110011011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111110000011010010011101010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110001101000101001011110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111111001000110011000010100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111011100001110001100011101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111101100010110010111000100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110101011000111100101111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111110110010000010111011101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111101000110000001100000010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111110011010011000110111000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111100100001000111110111011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111101101101110100001001100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111101101000111101000101110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111100100110010010010100101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111111100101000011110010010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111100111100100110111110011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111101000010110011011011000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel31_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel31 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111110101100011010010101101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel31[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel31_Valid_Out)
	);
	Adder_32input add_k31(
		.Data1(Data_Out_Kernel31[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel31[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel31[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel31[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel31[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel31[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel31[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel31[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel31[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel31[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel31[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel31[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel31[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel31[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel31[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel31[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel31[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel31[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel31[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel31[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel31[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel31[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel31[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel31[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel31[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel31[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel31[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel31[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel31[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel31[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel31[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel31[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel31),
		.Data_Out(add_k31_Data_Out),
		.Valid_Out(add_kernel31_Valid_Out)
	);
	Batch_Norm bn_kernel31(
		.Data_A(32'b00111110010011111100101110000100),
		.Data_B(32'b00111111100001100011110101010111),
		.Data_In(add_k31_Data_Out),
		.Valid_In(add_kernel31_Valid_Out),
		.Data_Out(bn31_Data_Out),
		.Valid_Out(bn31_Valid_Out)
	);
	Relu_Core rl_kernel31(
		.Data_In(bn31_Data_Out),
		.Valid_In(bn31_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(rl31_Valid_Out)
	);
//////////KERNEL32//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111110111001100010001011101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111101011110100110100011000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111100110000111101011011110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110110010101001100110110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111110101000100001110000001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110111001010010100100011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111110100000101010011111111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111110110100100100011110111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111101010001010100110111010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111110100100001001010111000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111110101011000011010001111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111111001110010000000000011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111100101100100000100000000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111111000100110010001000100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111101110001110111110111011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111101011100011010001000111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111111011000011110101111101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110001100100011110111101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111101100010010101100000111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111111000011110100010111010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110001000010000101010001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111110101010000011110111001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111110111011111001110111111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111110111010110100000011001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111110000100001111000000011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111110101101110100001110001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110111101100000001001111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111110010010101111101110101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111101110101010011001111001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111110110110100111101110110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111011101010011101111101000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel32_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel32 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111110000101011011001110110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel32[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel32_Valid_Out)
	);
	Adder_32input add_k32(
		.Data1(Data_Out_Kernel32[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel32[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel32[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel32[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel32[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel32[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel32[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel32[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel32[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel32[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel32[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel32[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel32[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel32[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel32[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel32[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel32[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel32[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel32[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel32[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel32[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel32[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel32[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel32[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel32[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel32[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel32[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel32[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel32[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel32[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel32[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel32[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel32),
		.Data_Out(add_k32_Data_Out),
		.Valid_Out(add_kernel32_Valid_Out)
	);
	Batch_Norm bn_kernel32(
		.Data_A(32'b00111110100000111111010111100110),
		.Data_B(32'b10111110100001000010010111011110),
		.Data_In(add_k32_Data_Out),
		.Valid_In(add_kernel32_Valid_Out),
		.Data_Out(bn32_Data_Out),
		.Valid_Out(bn32_Valid_Out)
	);
	Relu_Core rl_kernel32(
		.Data_In(bn32_Data_Out),
		.Valid_In(bn32_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(rl32_Valid_Out)
	);
//////////KERNEL33//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110011000000001000001100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111110111011011110001010001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110010010100000101011110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111101100100101001101110110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111111010011101100111001101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111101101000011101010100010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111111011101111111101000111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111110010101010001000000001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111111000100100000001010010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111110000001001111011110010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110001001010101111010011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110100001001001010101011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110101100100011000111000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111110010101010101010111101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111101110101010011010100001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111110111100001101111001110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110000111111101001101001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110111001101111110001010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110011000000010100010001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110100001001110110100111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111101101111000101000010101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111110111110100100100100001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111110110100011010001101110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111110110001111000000100001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111101101110111111001001101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111111000100101011001111111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110111001000011100111110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110000001110110111011011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111110101000100011101001011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111100101111000111111000000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111110100011001111011111111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel33_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel33 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110110000010000001011100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel33[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel33_Valid_Out)
	);
	Adder_32input add_k33(
		.Data1(Data_Out_Kernel33[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel33[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel33[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel33[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel33[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel33[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel33[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel33[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel33[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel33[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel33[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel33[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel33[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel33[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel33[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel33[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel33[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel33[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel33[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel33[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel33[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel33[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel33[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel33[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel33[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel33[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel33[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel33[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel33[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel33[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel33[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel33[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel33),
		.Data_Out(add_k33_Data_Out),
		.Valid_Out(add_kernel33_Valid_Out)
	);
	Batch_Norm bn_kernel33(
		.Data_A(32'b00111110011011101000001011101000),
		.Data_B(32'b00111110100000001001100001011010),
		.Data_In(add_k33_Data_Out),
		.Valid_In(add_kernel33_Valid_Out),
		.Data_Out(bn33_Data_Out),
		.Valid_Out(bn33_Valid_Out)
	);
	Relu_Core rl_kernel33(
		.Data_In(bn33_Data_Out),
		.Valid_In(bn33_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*33-1:DATA_WIDHT*32]),
		.Valid_Out(rl33_Valid_Out)
	);
//////////KERNEL34//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111110100110110110010001101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111100111010110001100010101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111011101100000000000111101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111100001001000100111110110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111110100111001010011110000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111110000100010011110100100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111110100111100010001010101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111110110110111101100000100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110100110001110110101011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111110000100111110010010011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111110111100101010010100100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111110100101100111010011000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111101110001111011110010010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111110001100111101010111001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110100110011101110010000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111110100010100110010111100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111110000001000100110011011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111111000111100111011000000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111110110110001101101000001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111101111011101001000010100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110101111010100011010101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111110101111001111010111101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111110010011001111001101011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111100010000101000101100110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111110010010110010000101110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110001000000011111101101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111110110000110101101000110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111111001111000010011100100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111110101110110101100010000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111101001011111101111011000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111111011100111100001100100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel34_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel34 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111111001000010101100111110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel34[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel34_Valid_Out)
	);
	Adder_32input add_k34(
		.Data1(Data_Out_Kernel34[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel34[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel34[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel34[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel34[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel34[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel34[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel34[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel34[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel34[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel34[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel34[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel34[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel34[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel34[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel34[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel34[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel34[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel34[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel34[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel34[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel34[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel34[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel34[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel34[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel34[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel34[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel34[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel34[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel34[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel34[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel34[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel34),
		.Data_Out(add_k34_Data_Out),
		.Valid_Out(add_kernel34_Valid_Out)
	);
	Batch_Norm bn_kernel34(
		.Data_A(32'b00111110011010110100001110010101),
		.Data_B(32'b00111101101000100001001011111001),
		.Data_In(add_k34_Data_Out),
		.Valid_In(add_kernel34_Valid_Out),
		.Data_Out(bn34_Data_Out),
		.Valid_Out(bn34_Valid_Out)
	);
	Relu_Core rl_kernel34(
		.Data_In(bn34_Data_Out),
		.Valid_In(bn34_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*34-1:DATA_WIDHT*33]),
		.Valid_Out(rl34_Valid_Out)
	);
//////////KERNEL35//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111101101100010001001010101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111101110110110100010001011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111101011010111101100010011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110010111111010100011010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111111001011101000100101100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111101000111101001110111101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111110100110011111000010010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111110001001111000110111101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111110101000000010101101010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111110100100001101111100010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110111101000101011110001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111111000010001000000111011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111110011110000101011101110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111111000100111101011011000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110111111011010100011000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111110100110101101000110100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111100110010111010001000111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110100100100110101111111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111101011100001000110010111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111101110000010000011011101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110010110110100000000010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111110010000000011110010110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111111100101001010011111000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111110011101100000110010010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111110001011010000010110111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110001011100111001010001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110010000111000011000001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110101010100011011101110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111110101001000111000000000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111110110111111001101011001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111110100010011001111010001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel35_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel35 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111110110011111010101001000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel35[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel35_Valid_Out)
	);
	Adder_32input add_k35(
		.Data1(Data_Out_Kernel35[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel35[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel35[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel35[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel35[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel35[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel35[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel35[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel35[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel35[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel35[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel35[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel35[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel35[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel35[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel35[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel35[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel35[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel35[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel35[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel35[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel35[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel35[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel35[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel35[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel35[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel35[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel35[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel35[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel35[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel35[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel35[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel35),
		.Data_Out(add_k35_Data_Out),
		.Valid_Out(add_kernel35_Valid_Out)
	);
	Batch_Norm bn_kernel35(
		.Data_A(32'b00111110011010010011100100011000),
		.Data_B(32'b10111011011001011110000101100100),
		.Data_In(add_k35_Data_Out),
		.Valid_In(add_kernel35_Valid_Out),
		.Data_Out(bn35_Data_Out),
		.Valid_Out(bn35_Valid_Out)
	);
	Relu_Core rl_kernel35(
		.Data_In(bn35_Data_Out),
		.Valid_In(bn35_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*35-1:DATA_WIDHT*34]),
		.Valid_Out(rl35_Valid_Out)
	);
//////////KERNEL36//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111111001100111001010011000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111111011110011111111111001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110000000111110001101100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110110011010111111010101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111110110100111000011110010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111110100110011101000001111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111110001010111110100001110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111101010111001010100000101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111111000101110000111011001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111110001111111000000110000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111110110001011101001010111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111110011101010100001001100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111111010010001101011111011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111110011011001101111011100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110001011001110001100011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111110010101101011010011011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111110001101011111000111001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111110010110100100000000010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110111111011001010010101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111110011010111000000011110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111101110101111000110010110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111110010110001000010111011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111110111011111001100110010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111110110011100000101101011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111110000110010010100101000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111111000100011100101111000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111101100110111010010001100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110011111001111110000101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111101000101011000011111100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111110001110001110110000011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111110101110101001010001001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel36_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel36 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110100111111101011101001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel36[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel36_Valid_Out)
	);
	Adder_32input add_k36(
		.Data1(Data_Out_Kernel36[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel36[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel36[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel36[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel36[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel36[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel36[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel36[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel36[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel36[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel36[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel36[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel36[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel36[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel36[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel36[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel36[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel36[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel36[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel36[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel36[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel36[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel36[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel36[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel36[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel36[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel36[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel36[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel36[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel36[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel36[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel36[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel36),
		.Data_Out(add_k36_Data_Out),
		.Valid_Out(add_kernel36_Valid_Out)
	);
	Batch_Norm bn_kernel36(
		.Data_A(32'b00111110011101011010000000001010),
		.Data_B(32'b10111101101101100001011011010101),
		.Data_In(add_k36_Data_Out),
		.Valid_In(add_kernel36_Valid_Out),
		.Data_Out(bn36_Data_Out),
		.Valid_Out(bn36_Valid_Out)
	);
	Relu_Core rl_kernel36(
		.Data_In(bn36_Data_Out),
		.Valid_In(bn36_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*36-1:DATA_WIDHT*35]),
		.Valid_Out(rl36_Valid_Out)
	);
//////////KERNEL37//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111110101010011100100011100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111100111001001010001001000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110101001010011010110001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111100111101011111110101110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111110100000110001000010101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111011100000111010001101101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111111010000010011001001100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111110101000111100101010000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110100111011101100001011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111111000010101111001001111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111111000000010110101111010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110001100111110001000001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110100100011001001100110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111110110111101011001001000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110011110110011111110001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111110010010001101010010110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111111001011011111111100111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111110111010110011100001000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110100111101100101111100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110101110110011100100011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110010001100110010100100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111110111101111110001101011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111001011100001111010000111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111110110001110100010111101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111110100011001010011101011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111101100011100100101110100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111110011000110000000010100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111011110110011100000001100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111110101101101010001000000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111110001101111000100101101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111111010101100110100111110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel37_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel37 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111110010000100000000100010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel37[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel37_Valid_Out)
	);
	Adder_32input add_k37(
		.Data1(Data_Out_Kernel37[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel37[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel37[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel37[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel37[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel37[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel37[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel37[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel37[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel37[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel37[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel37[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel37[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel37[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel37[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel37[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel37[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel37[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel37[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel37[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel37[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel37[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel37[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel37[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel37[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel37[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel37[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel37[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel37[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel37[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel37[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel37[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel37),
		.Data_Out(add_k37_Data_Out),
		.Valid_Out(add_kernel37_Valid_Out)
	);
	Batch_Norm bn_kernel37(
		.Data_A(32'b00111110011101111001001110100001),
		.Data_B(32'b00111110010011010001010011010111),
		.Data_In(add_k37_Data_Out),
		.Valid_In(add_kernel37_Valid_Out),
		.Data_Out(bn37_Data_Out),
		.Valid_Out(bn37_Valid_Out)
	);
	Relu_Core rl_kernel37(
		.Data_In(bn37_Data_Out),
		.Valid_In(bn37_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*37-1:DATA_WIDHT*36]),
		.Valid_Out(rl37_Valid_Out)
	);
//////////KERNEL38//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111101100110001100110110110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110101010000101010110011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110101001010101000011010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110110001101001100101100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111110110101100100101010110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110111110101110111101100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111110100100000101100011011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111011110000000101110111110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111110110010011111010000111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111110111010110001011111111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110001101001101111101001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110101000100010011100111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111101100001110010111110111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111101010100110101110111100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110000110111111110011011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111111010000100100100101110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111110111000000010111101011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110001100110101100010110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111100100000101101111101100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111111010010100111010010001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111111010001101101000000110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111110110001001111111101101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111110101110100011010010001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111110100011110100001101000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111110001111001000100000111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111110110000101001111110011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111110100011110001000111100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111110101101010000011110100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111110110101011110100010000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111110101010101101010011100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111110100111011110001011101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel38_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel38 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111110110100100101000000100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel38[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel38_Valid_Out)
	);
	Adder_32input add_k38(
		.Data1(Data_Out_Kernel38[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel38[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel38[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel38[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel38[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel38[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel38[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel38[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel38[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel38[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel38[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel38[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel38[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel38[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel38[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel38[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel38[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel38[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel38[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel38[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel38[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel38[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel38[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel38[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel38[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel38[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel38[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel38[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel38[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel38[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel38[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel38[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel38),
		.Data_Out(add_k38_Data_Out),
		.Valid_Out(add_kernel38_Valid_Out)
	);
	Batch_Norm bn_kernel38(
		.Data_A(32'b00111110100000001111000110000011),
		.Data_B(32'b00111111010111100110000011100000),
		.Data_In(add_k38_Data_Out),
		.Valid_In(add_kernel38_Valid_Out),
		.Data_Out(bn38_Data_Out),
		.Valid_Out(bn38_Valid_Out)
	);
	Relu_Core rl_kernel38(
		.Data_In(bn38_Data_Out),
		.Valid_In(bn38_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*38-1:DATA_WIDHT*37]),
		.Valid_Out(rl38_Valid_Out)
	);
//////////KERNEL39//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111110110001001010101101111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111111000101111110110110111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111101111011100000101000110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110110010011010011100100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111110000110100010000111111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111110100010110001001110001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111110111010100110001111011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111100110011000010011001111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110101101101010000110110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111101110001111110010111110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110100001000010100100000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111110100100010111011000111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111111000101010110100010000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111110110111110111010001100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110100101000000011101010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111110010111101011000011111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110111001110001111100000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111110100010011101000111101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111101100000101110110011000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111110110100001100010010010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111100001110101001111101111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111110001110000110010011000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111111000010101101100101000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111111000001110111011011110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111110101110010100001111101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111110110010010000111010101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111110111100011010100000010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111111011011011111100101111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111110100111001001111011110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111101011100101000001010101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111110100111001110110110000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel39_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel39 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111101100000110011000100010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel39[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel39_Valid_Out)
	);
	Adder_32input add_k39(
		.Data1(Data_Out_Kernel39[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel39[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel39[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel39[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel39[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel39[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel39[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel39[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel39[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel39[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel39[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel39[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel39[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel39[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel39[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel39[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel39[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel39[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel39[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel39[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel39[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel39[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel39[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel39[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel39[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel39[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel39[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel39[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel39[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel39[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel39[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel39[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel39),
		.Data_Out(add_k39_Data_Out),
		.Valid_Out(add_kernel39_Valid_Out)
	);
	Batch_Norm bn_kernel39(
		.Data_A(32'b00111110100001010010111011000011),
		.Data_B(32'b10111111100111001111010001011101),
		.Data_In(add_k39_Data_Out),
		.Valid_In(add_kernel39_Valid_Out),
		.Data_Out(bn39_Data_Out),
		.Valid_Out(bn39_Valid_Out)
	);
	Relu_Core rl_kernel39(
		.Data_In(bn39_Data_Out),
		.Valid_In(bn39_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*39-1:DATA_WIDHT*38]),
		.Valid_Out(rl39_Valid_Out)
	);
//////////KERNEL40//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111110101000000101110010011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110110100100101100110101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111101001111011010101001010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111111010000110000001011001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111110001111100011111010111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111110000101011011111110011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111101101000000000001010010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111100000010001100111111010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110111000000010100010010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111101100011111111000000010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111111100000101000011100100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110111000111101001001010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111110001010111111011000100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111110100100010100110110001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110100100111101100011111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111110100111110100100001000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111101110101101001010010001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111110100010111110000001101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110001110111010001111011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111101110011010101110011100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110000000100011111101110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111111000100011000111101010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110111000011110110011000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111111001111011000111110111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111110001101101100101101001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111101100001010111010010011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111110011100111000111011001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111110010101101001010111000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111100101100101110001010111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111110101101011111010111010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111111001001111001010110111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel40_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel40 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111101101001001100110111010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel40[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel40_Valid_Out)
	);
	Adder_32input add_k40(
		.Data1(Data_Out_Kernel40[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel40[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel40[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel40[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel40[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel40[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel40[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel40[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel40[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel40[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel40[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel40[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel40[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel40[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel40[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel40[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel40[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel40[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel40[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel40[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel40[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel40[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel40[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel40[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel40[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel40[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel40[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel40[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel40[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel40[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel40[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel40[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel40),
		.Data_Out(add_k40_Data_Out),
		.Valid_Out(add_kernel40_Valid_Out)
	);
	Batch_Norm bn_kernel40(
		.Data_A(32'b00111110011111110000011000000000),
		.Data_B(32'b00111110111111010011001101101111),
		.Data_In(add_k40_Data_Out),
		.Valid_In(add_kernel40_Valid_Out),
		.Data_Out(bn40_Data_Out),
		.Valid_Out(bn40_Valid_Out)
	);
	Relu_Core rl_kernel40(
		.Data_In(bn40_Data_Out),
		.Valid_In(bn40_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*40-1:DATA_WIDHT*39]),
		.Valid_Out(rl40_Valid_Out)
	);
//////////KERNEL41//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111110100001111101101111111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111101101010100010000111011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110111110010010001011000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111101111011110011011010000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111111000111111100010100110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111110100101010001111000011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111110010110110011101011010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111110011101001010001010000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111101100011010011011110010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111111010101101111000001110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111101001101000101111100101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111110010011110110111110000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110010010100110100010110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111101000001111010000111101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111101011100101000011110011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111110100000111000011001011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111101100111100011000110111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111110111101110101001101001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111111000110001001100111011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110110100101000111001100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110110110000001110011100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111111000111100011100111011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110100110000010101000001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111101100011011000010101001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111110101000101010110000101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111011111100110011000110001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111100100101111001111011101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111111001001111001001111001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111101010100000110101011111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110111111111011011100000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111111000010100110011110100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel41_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel41 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111111000010100011011101010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel41[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel41_Valid_Out)
	);
	Adder_32input add_k41(
		.Data1(Data_Out_Kernel41[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel41[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel41[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel41[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel41[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel41[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel41[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel41[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel41[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel41[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel41[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel41[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel41[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel41[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel41[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel41[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel41[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel41[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel41[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel41[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel41[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel41[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel41[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel41[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel41[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel41[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel41[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel41[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel41[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel41[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel41[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel41[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel41),
		.Data_Out(add_k41_Data_Out),
		.Valid_Out(add_kernel41_Valid_Out)
	);
	Batch_Norm bn_kernel41(
		.Data_A(32'b00111110100001100100001101000101),
		.Data_B(32'b00111110011101111011111110100100),
		.Data_In(add_k41_Data_Out),
		.Valid_In(add_kernel41_Valid_Out),
		.Data_Out(bn41_Data_Out),
		.Valid_Out(bn41_Valid_Out)
	);
	Relu_Core rl_kernel41(
		.Data_In(bn41_Data_Out),
		.Valid_In(bn41_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*41-1:DATA_WIDHT*40]),
		.Valid_Out(rl41_Valid_Out)
	);
//////////KERNEL42//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111111001011000100001010101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111101110101101100001111100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111111001101100100000101010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110011101110101101001011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111110001011001101101110111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111111001110011010001110011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111110001100000011001000110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111110101100001000111000110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111111000001100000100110001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111110010101100110101010111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111110101011010101100100110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110011100011001001111100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111110100111100101001101000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111110101001111100001001100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110010001000100010001000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111101100101100010101011101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111111010110111000110110011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111110110111111010101101111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111110110110110100100110000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111011000110001001111110110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110011011000110010101101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111110011100110000000101110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111110011100000101001111010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111101001001000011010011100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111101111010001011111101001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111110011101100011011000111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111111000100000010011000110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111011101010111011010111100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111101000010101110110111001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111101111100000101100111011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111110100100010101110000101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel42_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel42 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111110101111110010010011011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel42[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel42_Valid_Out)
	);
	Adder_32input add_k42(
		.Data1(Data_Out_Kernel42[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel42[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel42[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel42[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel42[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel42[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel42[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel42[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel42[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel42[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel42[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel42[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel42[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel42[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel42[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel42[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel42[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel42[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel42[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel42[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel42[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel42[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel42[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel42[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel42[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel42[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel42[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel42[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel42[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel42[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel42[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel42[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel42),
		.Data_Out(add_k42_Data_Out),
		.Valid_Out(add_kernel42_Valid_Out)
	);
	Batch_Norm bn_kernel42(
		.Data_A(32'b00111110010111110100111001111101),
		.Data_B(32'b10111100111111111100100110110011),
		.Data_In(add_k42_Data_Out),
		.Valid_In(add_kernel42_Valid_Out),
		.Data_Out(bn42_Data_Out),
		.Valid_Out(bn42_Valid_Out)
	);
	Relu_Core rl_kernel42(
		.Data_In(bn42_Data_Out),
		.Valid_In(bn42_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*42-1:DATA_WIDHT*41]),
		.Valid_Out(rl42_Valid_Out)
	);
//////////KERNEL43//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110101001100110011100010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110110001001111110101000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111101010011011000110001101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110100001011010001101000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111111100010011100110111101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111110010010000111010010001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111101100000110011111101011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111110110010111010101111000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111110000101110010001110010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111101100100100110000111001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111100100100100100001010011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111110110001101010101000110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111101010001100000000110011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111110001010010011010001101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110010000101100011000101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111110100010101111010011111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111111000110000011001001101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111111000101100010111011001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111100100011100111100011100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110100010111101100010011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110111100110001111101110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111110000100101001101000100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111100110111000111010011000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111110000101011011111101010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111111000110011101011100011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111110010000100001011101001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110011000010110101101100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111101011000100100000100101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111110110011111111000011110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111111010000101110101110001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111110110011010101110101000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel43_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel43 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111110010011100110001101101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel43[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel43_Valid_Out)
	);
	Adder_32input add_k43(
		.Data1(Data_Out_Kernel43[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel43[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel43[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel43[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel43[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel43[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel43[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel43[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel43[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel43[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel43[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel43[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel43[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel43[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel43[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel43[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel43[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel43[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel43[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel43[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel43[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel43[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel43[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel43[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel43[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel43[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel43[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel43[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel43[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel43[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel43[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel43[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel43),
		.Data_Out(add_k43_Data_Out),
		.Valid_Out(add_kernel43_Valid_Out)
	);
	Batch_Norm bn_kernel43(
		.Data_A(32'b00111110100101110001010101010001),
		.Data_B(32'b10111110010011110010000100111110),
		.Data_In(add_k43_Data_Out),
		.Valid_In(add_kernel43_Valid_Out),
		.Data_Out(bn43_Data_Out),
		.Valid_Out(bn43_Valid_Out)
	);
	Relu_Core rl_kernel43(
		.Data_In(bn43_Data_Out),
		.Valid_In(bn43_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*43-1:DATA_WIDHT*42]),
		.Valid_Out(rl43_Valid_Out)
	);
//////////KERNEL44//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111110100100010001001011011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111110010000100001011110010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110011111001011110000101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110101110010011000000101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111011101111100110001110011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111110110001101101001011000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111110000010101100011101010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111110001111111100010000010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110011001111101101010110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111111001000100010101011110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111100111111010111110010010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111110110000000010111001101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110110101111111101010100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111100011110001010110011011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111111010101110111101011011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111111000011011000000001111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111110000011111011100001010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110010100001111010100111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111100001010010010010100000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111111010000100001011001110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110110000110011110001011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111101111111110110111001011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111110011101000010100100110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111110001111100100111101001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111111000010001100000000001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111110101011010110000100011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111110101010000110010000100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111110110010100011010111001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111100110100111110010000110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111101011000001011111110101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111111010000010111111101011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel44_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel44 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110100110111001100100110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel44[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel44_Valid_Out)
	);
	Adder_32input add_k44(
		.Data1(Data_Out_Kernel44[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel44[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel44[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel44[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel44[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel44[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel44[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel44[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel44[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel44[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel44[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel44[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel44[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel44[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel44[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel44[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel44[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel44[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel44[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel44[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel44[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel44[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel44[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel44[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel44[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel44[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel44[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel44[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel44[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel44[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel44[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel44[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel44),
		.Data_Out(add_k44_Data_Out),
		.Valid_Out(add_kernel44_Valid_Out)
	);
	Batch_Norm bn_kernel44(
		.Data_A(32'b00111110100100100100011100000011),
		.Data_B(32'b00111111010000100101001100010000),
		.Data_In(add_k44_Data_Out),
		.Valid_In(add_kernel44_Valid_Out),
		.Data_Out(bn44_Data_Out),
		.Valid_Out(bn44_Valid_Out)
	);
	Relu_Core rl_kernel44(
		.Data_In(bn44_Data_Out),
		.Valid_In(bn44_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*44-1:DATA_WIDHT*43]),
		.Valid_Out(rl44_Valid_Out)
	);
//////////KERNEL45//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111111001001001110010110110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110011100110001110001011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111111000111101101000101111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110100011110100001010010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111110010110011110111100101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111101100100101000101101001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111110010110101001111111011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111111001001011111010110010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111100100001011101110100011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110110101001100001110000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111110110010011111011011000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111101101001001100100000010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111101001111000001101111000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111110101000000100101000000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110001111111110110101100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111101101110101000111101100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110000101000010000100011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111110101000010101000011011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111110111111111000111110011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111111001100011110110011010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110000110101000101100010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111110111110111000110111100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111111000100000011000000101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111111010000101000000110101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111110111110101000101010100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111101000011011000010111100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111100110101100000100101000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110011111010011011011000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111111000010101000011110000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111101100011010110000111000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111101100100000111101000111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel45_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel45 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111101111111110111110001110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel45[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel45_Valid_Out)
	);
	Adder_32input add_k45(
		.Data1(Data_Out_Kernel45[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel45[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel45[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel45[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel45[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel45[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel45[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel45[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel45[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel45[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel45[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel45[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel45[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel45[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel45[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel45[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel45[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel45[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel45[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel45[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel45[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel45[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel45[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel45[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel45[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel45[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel45[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel45[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel45[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel45[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel45[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel45[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel45),
		.Data_Out(add_k45_Data_Out),
		.Valid_Out(add_kernel45_Valid_Out)
	);
	Batch_Norm bn_kernel45(
		.Data_A(32'b00111110010011100111001011011011),
		.Data_B(32'b10111111100000111011111100011001),
		.Data_In(add_k45_Data_Out),
		.Valid_In(add_kernel45_Valid_Out),
		.Data_Out(bn45_Data_Out),
		.Valid_Out(bn45_Valid_Out)
	);
	Relu_Core rl_kernel45(
		.Data_In(bn45_Data_Out),
		.Valid_In(bn45_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*45-1:DATA_WIDHT*44]),
		.Valid_Out(rl45_Valid_Out)
	);
//////////KERNEL46//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111110101010010100010111110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110100110110001001111010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110111010100110100100001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110010110010110010011101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111110101010010011010101111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111110100010000001000001110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111101101000011110111001001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111110000000100100000110000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111110010011100110110101010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111110000111110011000010000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111110000010110010011000101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111101011001110101111010011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111101010100001110010100000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111110110101011110010001001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111111000110100011111010110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111110101001010011001000100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110101110001101111010110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110100001010001000111010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111111010111110101100101011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111110011110001001101011011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110101000100000101010110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111101000110110111110110111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111111000011000011010111010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111110110101110100110111000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111110000110000100001001001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110110111110001011000110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110011101111111111011000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111111000010011111001010101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111110010011110000001110011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111111000010001011011100011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111110000110100101100100100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel46_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel46 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111111010011110001011010000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel46[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel46_Valid_Out)
	);
	Adder_32input add_k46(
		.Data1(Data_Out_Kernel46[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel46[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel46[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel46[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel46[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel46[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel46[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel46[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel46[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel46[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel46[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel46[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel46[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel46[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel46[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel46[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel46[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel46[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel46[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel46[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel46[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel46[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel46[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel46[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel46[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel46[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel46[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel46[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel46[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel46[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel46[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel46[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel46),
		.Data_Out(add_k46_Data_Out),
		.Valid_Out(add_kernel46_Valid_Out)
	);
	Batch_Norm bn_kernel46(
		.Data_A(32'b00111110100011011110000000000011),
		.Data_B(32'b00111110000100100001010100100110),
		.Data_In(add_k46_Data_Out),
		.Valid_In(add_kernel46_Valid_Out),
		.Data_Out(bn46_Data_Out),
		.Valid_Out(bn46_Valid_Out)
	);
	Relu_Core rl_kernel46(
		.Data_In(bn46_Data_Out),
		.Valid_In(bn46_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*46-1:DATA_WIDHT*45]),
		.Valid_Out(rl46_Valid_Out)
	);
//////////KERNEL47//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111111000110110100110111100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110100000111110111110000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110101101100111011101100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110100101110101100110100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111101001110101111100101000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111101110101110101000110100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111101111011110111100100100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111101011111111101100010011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110111111010110111100000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110110001011001110101001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110100110011001110001000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111101010101011111100100011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111100111111111101001001010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111111001010100110001000001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110101110000000010011000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111110100001010100110010001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111110111010110110000111101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111101100011101111101110100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110110001110111100000000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110100110010010100100100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110001001110111110001101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111101001101111010000001110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111101110110100000001011011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111101100001111000001110110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111101010100111100101010010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111111001011000111101011000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110101100111101001001100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110111100111000000011001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111110001011111010111101001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111101100000100000011101111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111111001101011011010100101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel47_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel47 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111111000111011111001010101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel47[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel47_Valid_Out)
	);
	Adder_32input add_k47(
		.Data1(Data_Out_Kernel47[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel47[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel47[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel47[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel47[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel47[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel47[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel47[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel47[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel47[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel47[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel47[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel47[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel47[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel47[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel47[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel47[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel47[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel47[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel47[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel47[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel47[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel47[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel47[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel47[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel47[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel47[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel47[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel47[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel47[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel47[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel47[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel47),
		.Data_Out(add_k47_Data_Out),
		.Valid_Out(add_kernel47_Valid_Out)
	);
	Batch_Norm bn_kernel47(
		.Data_A(32'b00111110100011100000000101010010),
		.Data_B(32'b10111111100011000100011110110100),
		.Data_In(add_k47_Data_Out),
		.Valid_In(add_kernel47_Valid_Out),
		.Data_Out(bn47_Data_Out),
		.Valid_Out(bn47_Valid_Out)
	);
	Relu_Core rl_kernel47(
		.Data_In(bn47_Data_Out),
		.Valid_In(bn47_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*47-1:DATA_WIDHT*46]),
		.Valid_Out(rl47_Valid_Out)
	);
//////////KERNEL48//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111110111011110011001100111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111110110010010101111101000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111111000111100011010000100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110011111000111100001001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111110000111100011010001011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110111000110011111010100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111110000001111100110110001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111110101010000010100111010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111111001100010010010001010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111111001000011110110011111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111101101010011101011011010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110100001111001100000000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111110001001111110011000110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111110110001100011111011001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110110010110011000101101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111111001101011110100011100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111111001111111100011010100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110101101100100101000100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111110011000011100110110011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111110011011110100110011010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111101100000111000011101000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111101101110011101101000011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110010110101101011010011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111110110001100110001101010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111110010010100010001101000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110011001011111010110110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111101101111011110011001101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110011001101010000110110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111110011001010100111010000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110000111001011010001001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111110101011100110001011011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel48_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel48 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111110000001001111010011000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel48[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel48_Valid_Out)
	);
	Adder_32input add_k48(
		.Data1(Data_Out_Kernel48[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel48[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel48[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel48[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel48[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel48[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel48[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel48[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel48[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel48[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel48[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel48[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel48[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel48[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel48[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel48[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel48[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel48[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel48[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel48[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel48[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel48[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel48[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel48[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel48[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel48[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel48[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel48[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel48[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel48[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel48[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel48[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel48),
		.Data_Out(add_k48_Data_Out),
		.Valid_Out(add_kernel48_Valid_Out)
	);
	Batch_Norm bn_kernel48(
		.Data_A(32'b00111110011111010011000000111010),
		.Data_B(32'b00111110100110100001001000100100),
		.Data_In(add_k48_Data_Out),
		.Valid_In(add_kernel48_Valid_Out),
		.Data_Out(bn48_Data_Out),
		.Valid_Out(bn48_Valid_Out)
	);
	Relu_Core rl_kernel48(
		.Data_In(bn48_Data_Out),
		.Valid_In(bn48_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*48-1:DATA_WIDHT*47]),
		.Valid_Out(rl48_Valid_Out)
	);
//////////KERNEL49//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111101110000111110100100111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111101110100101110001111001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110100000001111110000100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110100111111010101100000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111101100000000100110001111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111110010000111011010001011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111111001111000100010000011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111110100000110100110000010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111110011010101100011010111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111101101100000100100111101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110011111011011001111010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111110110100101010010101010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110101101011001001001111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111110100100111111100110110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111101000001011100010000000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111110101101001001001101010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111111010011001010100011010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110001100110001001101101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110110001011001011001101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111110110101110011101010101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111111000010010111011000100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111101100000100001100111110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111110100000110001110100101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111110110010000011110111001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111101011000011101100001011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111100010100111010011111111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111101110111011100101110111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111111000001000111010100000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111111011101110001010000001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110110000000010010100100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111101000010110011110110111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel49_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel49 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110001100000011111000001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel49[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel49_Valid_Out)
	);
	Adder_32input add_k49(
		.Data1(Data_Out_Kernel49[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel49[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel49[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel49[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel49[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel49[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel49[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel49[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel49[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel49[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel49[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel49[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel49[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel49[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel49[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel49[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel49[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel49[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel49[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel49[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel49[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel49[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel49[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel49[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel49[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel49[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel49[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel49[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel49[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel49[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel49[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel49[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel49),
		.Data_Out(add_k49_Data_Out),
		.Valid_Out(add_kernel49_Valid_Out)
	);
	Batch_Norm bn_kernel49(
		.Data_A(32'b00111110010101100000101010100101),
		.Data_B(32'b00111101100101110110110111001101),
		.Data_In(add_k49_Data_Out),
		.Valid_In(add_kernel49_Valid_Out),
		.Data_Out(bn49_Data_Out),
		.Valid_Out(bn49_Valid_Out)
	);
	Relu_Core rl_kernel49(
		.Data_In(bn49_Data_Out),
		.Valid_In(bn49_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*49-1:DATA_WIDHT*48]),
		.Valid_Out(rl49_Valid_Out)
	);
//////////KERNEL50//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110100100110001101110010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110101010101110111001011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111111000010001000100110011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110011111001111011101011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111101100000011010111001110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111101001101010101000010000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111101011100001111101011011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111110000100101011001010011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110011111011101011111101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110100111001000111101001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111111000011101001100111011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111111001010100000101111010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110011100000111101011010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111110100111011011101010110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110111001010110011100000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111110100000010100100011010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111111000110100100001010101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110100100110010110000110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111111000011011001101010101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111111011110011010100011110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110000000111000111000111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111111010000001010101101001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111110001101101000010100010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111110001011101100101000010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111100110101101100110101000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111111001000011100101100100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110001001100111111111001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111100011010100111011010000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111101101001011001100010010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111101000111100101110100101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111101010110110101111101001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel50_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel50 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110100101101100011101001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel50[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel50_Valid_Out)
	);
	Adder_32input add_k50(
		.Data1(Data_Out_Kernel50[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel50[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel50[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel50[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel50[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel50[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel50[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel50[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel50[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel50[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel50[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel50[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel50[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel50[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel50[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel50[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel50[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel50[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel50[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel50[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel50[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel50[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel50[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel50[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel50[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel50[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel50[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel50[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel50[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel50[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel50[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel50[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel50),
		.Data_Out(add_k50_Data_Out),
		.Valid_Out(add_kernel50_Valid_Out)
	);
	Batch_Norm bn_kernel50(
		.Data_A(32'b00111110100010010110010110100001),
		.Data_B(32'b10111111100000000101010100101111),
		.Data_In(add_k50_Data_Out),
		.Valid_In(add_kernel50_Valid_Out),
		.Data_Out(bn50_Data_Out),
		.Valid_Out(bn50_Valid_Out)
	);
	Relu_Core rl_kernel50(
		.Data_In(bn50_Data_Out),
		.Valid_In(bn50_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*50-1:DATA_WIDHT*49]),
		.Valid_Out(rl50_Valid_Out)
	);
//////////KERNEL51//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110101110100101010010100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111011001110010100100111101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111100000110011111101001001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111111000011011100011000110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111111010010100100111110001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110011110101010001001101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111110111110010011001111100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111101001101110111011000000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111110011001101110111001011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111101101011011111101010001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111110001011001001011000010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111110010010011000100100000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111101010101001101001111101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111101110011100010010000010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110001011001101011100100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111111000010000111111000111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111111000100010111111110111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111110000001110101001101001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111101101000011111011100111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110000101010101111001000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110101011101011111110100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111110011010111001100100110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111110111010000110111100100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111110110100110100011010001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111110101011010111100000110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111010001100000010011111110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110111010000001001000011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110000111110100111101011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111110101101101001001101010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111110101110001011101001001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111110100001101011000110110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel51_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel51 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111111001110000111011100001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel51[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel51_Valid_Out)
	);
	Adder_32input add_k51(
		.Data1(Data_Out_Kernel51[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel51[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel51[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel51[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel51[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel51[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel51[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel51[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel51[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel51[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel51[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel51[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel51[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel51[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel51[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel51[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel51[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel51[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel51[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel51[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel51[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel51[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel51[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel51[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel51[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel51[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel51[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel51[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel51[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel51[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel51[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel51[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel51),
		.Data_Out(add_k51_Data_Out),
		.Valid_Out(add_kernel51_Valid_Out)
	);
	Batch_Norm bn_kernel51(
		.Data_A(32'b00111110011110101110001100011110),
		.Data_B(32'b10111111010001001110100100011101),
		.Data_In(add_k51_Data_Out),
		.Valid_In(add_kernel51_Valid_Out),
		.Data_Out(bn51_Data_Out),
		.Valid_Out(bn51_Valid_Out)
	);
	Relu_Core rl_kernel51(
		.Data_In(bn51_Data_Out),
		.Valid_In(bn51_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*51-1:DATA_WIDHT*50]),
		.Valid_Out(rl51_Valid_Out)
	);
//////////KERNEL52//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110000001001111000111110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110001101010001001001100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110101000101100000010100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110111011010111101100001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111101100100010001010011111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111111100001100000001010110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111110111010001001000011101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111110000110011011001111110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111111000011110110110101110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111101011101000000010101110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111110111000000101001001010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111110000110111110000110010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111110010100010100011000010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111011111100010011111101110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111110011111110101111100001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111111000100011010110110110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110001110001100011110010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111100101100100010100001110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111111000110100000000110100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110101011111111000111000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110111000111100000010010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111101101111111010011000110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111110110101111010000111011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111110011111000100010111111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111101111000010111100000011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110111101110101111100111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111110101000001101011111101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110001000000101000000110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111110001010010101101110010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111110100011000110110101101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111101011100101010011100100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel52_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel52 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110101011101001011011011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel52[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel52_Valid_Out)
	);
	Adder_32input add_k52(
		.Data1(Data_Out_Kernel52[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel52[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel52[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel52[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel52[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel52[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel52[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel52[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel52[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel52[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel52[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel52[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel52[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel52[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel52[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel52[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel52[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel52[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel52[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel52[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel52[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel52[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel52[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel52[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel52[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel52[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel52[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel52[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel52[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel52[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel52[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel52[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel52),
		.Data_Out(add_k52_Data_Out),
		.Valid_Out(add_kernel52_Valid_Out)
	);
	Batch_Norm bn_kernel52(
		.Data_A(32'b00111110011101101101000110010010),
		.Data_B(32'b10111111000110000001101010100111),
		.Data_In(add_k52_Data_Out),
		.Valid_In(add_kernel52_Valid_Out),
		.Data_Out(bn52_Data_Out),
		.Valid_Out(bn52_Valid_Out)
	);
	Relu_Core rl_kernel52(
		.Data_In(bn52_Data_Out),
		.Valid_In(bn52_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*52-1:DATA_WIDHT*51]),
		.Valid_Out(rl52_Valid_Out)
	);
//////////KERNEL53//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110100011010111001001010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111110000100001100110011001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111100110110101011110001000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110010000010000000010010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111110101110110011011001011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111100010111000010000000011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111110010100101011110100001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111110101110001010011110110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111110101100101111110010110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111101101100100111111110010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b00111110010101000101010011011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111101001001110100110010001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111110001011001101000101101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111110100000100010011011010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110100000101000110010000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111110001001001001100100000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110111001011000000000011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111100111011000101100011011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111111000001111100011111001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111110111110111010100111111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110001011000100100111000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111111010101010100001011010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111110010111001011100000101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111111010001100000000011110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111111011000010111000101101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111110110010110000001110000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111110111111111110011001000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111110010101001011001101110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111110010001101100101011001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111101110100011010100101101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111110111111001100000010010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel53_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel53 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110100111100011010101111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel53[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel53_Valid_Out)
	);
	Adder_32input add_k53(
		.Data1(Data_Out_Kernel53[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel53[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel53[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel53[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel53[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel53[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel53[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel53[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel53[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel53[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel53[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel53[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel53[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel53[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel53[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel53[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel53[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel53[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel53[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel53[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel53[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel53[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel53[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel53[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel53[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel53[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel53[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel53[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel53[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel53[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel53[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel53[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel53),
		.Data_Out(add_k53_Data_Out),
		.Valid_Out(add_kernel53_Valid_Out)
	);
	Batch_Norm bn_kernel53(
		.Data_A(32'b00111110100011010101110010100010),
		.Data_B(32'b10111101100101100011010111010000),
		.Data_In(add_k53_Data_Out),
		.Valid_In(add_kernel53_Valid_Out),
		.Data_Out(bn53_Data_Out),
		.Valid_Out(bn53_Valid_Out)
	);
	Relu_Core rl_kernel53(
		.Data_In(bn53_Data_Out),
		.Valid_In(bn53_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*53-1:DATA_WIDHT*52]),
		.Valid_Out(rl53_Valid_Out)
	);
//////////KERNEL54//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110110001100010101011100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111111000100101010111100000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111101110000111010100011011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110000101111111111110100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111110100001111001011011000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111110110010101110101110001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111111001100010011100010000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111101110011010000100011000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111110100111000111011110010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110001101110001101110001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111100000111100110011110000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111111000000110110100110010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110100011000000101101100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111110100011000000001010010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111111001010111011010000100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111110010111001111101000000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110101111010001101011000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111101010000101010111010001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111111001110101001101100101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111110111111000000101010010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110010010010000111110011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111110011011001001111011110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111110001001110101000101101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111110000001001010001011001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111110010000000010110010001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111110111100001010011011110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111101110011100010100000100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111111001111000011001111000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111110100010101111111001111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111101010101100111100100010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111110011010101011000100101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel54_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel54 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111110010111100011101011010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel54[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel54_Valid_Out)
	);
	Adder_32input add_k54(
		.Data1(Data_Out_Kernel54[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel54[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel54[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel54[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel54[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel54[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel54[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel54[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel54[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel54[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel54[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel54[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel54[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel54[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel54[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel54[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel54[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel54[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel54[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel54[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel54[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel54[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel54[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel54[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel54[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel54[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel54[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel54[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel54[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel54[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel54[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel54[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel54),
		.Data_Out(add_k54_Data_Out),
		.Valid_Out(add_kernel54_Valid_Out)
	);
	Batch_Norm bn_kernel54(
		.Data_A(32'b00111110100111111101110001100010),
		.Data_B(32'b10111110100100111111111001100011),
		.Data_In(add_k54_Data_Out),
		.Valid_In(add_kernel54_Valid_Out),
		.Data_Out(bn54_Data_Out),
		.Valid_Out(bn54_Valid_Out)
	);
	Relu_Core rl_kernel54(
		.Data_In(bn54_Data_Out),
		.Valid_In(bn54_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*54-1:DATA_WIDHT*53]),
		.Valid_Out(rl54_Valid_Out)
	);
//////////KERNEL55//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111111000000000100011111101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111110100110000100011001001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110010100000110001001001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111101111111001101001000010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111110010100001000101111110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111101101001011101111000000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111110100011100011011110111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111111001110001110111110001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110101111011110110000110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110111001111010111111100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111110111100100101011011111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111110101011100110010011101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111110100101000001111110111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111111000101100000101011011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111101001101000101001100001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111101100011010010010011000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111111001000100100010001010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111110111000000000000110011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111101001101010000011110001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111101100111011010100100011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110100100101100111000110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111110110001101100101001101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110101010101100101011110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111111001001100111010100100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111111000001100100111110100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111101111110110101011100110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111110100110111011011111011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111101101011100100010100111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111110100001100100101001010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111110001001001001110101001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111110100110010010110011110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel55_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel55 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111110111101100010001001010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel55[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel55_Valid_Out)
	);
	Adder_32input add_k55(
		.Data1(Data_Out_Kernel55[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel55[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel55[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel55[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel55[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel55[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel55[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel55[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel55[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel55[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel55[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel55[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel55[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel55[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel55[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel55[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel55[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel55[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel55[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel55[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel55[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel55[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel55[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel55[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel55[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel55[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel55[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel55[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel55[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel55[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel55[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel55[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel55),
		.Data_Out(add_k55_Data_Out),
		.Valid_Out(add_kernel55_Valid_Out)
	);
	Batch_Norm bn_kernel55(
		.Data_A(32'b00111110100000001010001001011101),
		.Data_B(32'b00111110001011101000011010010000),
		.Data_In(add_k55_Data_Out),
		.Valid_In(add_kernel55_Valid_Out),
		.Data_Out(bn55_Data_Out),
		.Valid_Out(bn55_Valid_Out)
	);
	Relu_Core rl_kernel55(
		.Data_In(bn55_Data_Out),
		.Valid_In(bn55_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*55-1:DATA_WIDHT*54]),
		.Valid_Out(rl55_Valid_Out)
	);
//////////KERNEL56//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111101011101111001101001000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110110111100010111101101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111110010100011100010111001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111101100010110000101010001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111110111101100001110000110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111101110000001101001011001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111110001101001101110111001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111110101100001000101100110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110011111000101011111111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111110100111011011010000111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111110100011100000001100001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111110111000011000101010000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110101000000100100001111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111110000101101010011010111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110100111101111101011110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111101010011111011010110001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111111010010000000001001100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110111011110010010100111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110111111100010111000011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111101101111111010111001010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110100011110010111101011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111110100001101110010001001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111111100000000000001000011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111110100010010111010110110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111110101101010100110111000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110010111101111100110010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111111000001111101001101101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111101110100001111111111011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111110101100110101010110010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111111010101001001110001110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111110100101000110010011111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel56_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel56 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111101100000001001110111100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel56[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel56_Valid_Out)
	);
	Adder_32input add_k56(
		.Data1(Data_Out_Kernel56[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel56[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel56[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel56[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel56[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel56[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel56[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel56[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel56[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel56[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel56[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel56[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel56[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel56[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel56[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel56[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel56[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel56[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel56[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel56[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel56[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel56[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel56[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel56[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel56[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel56[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel56[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel56[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel56[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel56[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel56[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel56[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel56),
		.Data_Out(add_k56_Data_Out),
		.Valid_Out(add_kernel56_Valid_Out)
	);
	Batch_Norm bn_kernel56(
		.Data_A(32'b00111110011111010000000111111000),
		.Data_B(32'b00111111100001000011100101000001),
		.Data_In(add_k56_Data_Out),
		.Valid_In(add_kernel56_Valid_Out),
		.Data_Out(bn56_Data_Out),
		.Valid_Out(bn56_Valid_Out)
	);
	Relu_Core rl_kernel56(
		.Data_In(bn56_Data_Out),
		.Valid_In(bn56_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*56-1:DATA_WIDHT*55]),
		.Valid_Out(rl56_Valid_Out)
	);
//////////KERNEL57//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111101100101001110000001101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110101000101101010111010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110100011101001001000100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110101100000000111101110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111110111100111010100110001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111111001001110100101010101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111110000100000111111001010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111101111111110110110100000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110101111100010110100101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111110011011011110010101111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111100111010000110000001011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111100110111010000101010111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110110011001100010011011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111100001111111111111010101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111101111001000000001110100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111110000111000000011011110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111110101001110010010111111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110010010000010111011110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111101101011111100001011011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111110001101011001001011110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111111001001101111110001011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111111000000010110101001000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111110101100100000101110000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111110100101010111000011011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111110101111011100001110000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111111010010000100100110100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111111011011111100101011010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111101100011100110100010011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111100011001011111011000110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111111010011110111100111101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111110010010010110100100010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel57_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel57 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b00111101111100010101110111000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel57[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel57_Valid_Out)
	);
	Adder_32input add_k57(
		.Data1(Data_Out_Kernel57[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel57[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel57[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel57[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel57[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel57[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel57[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel57[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel57[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel57[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel57[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel57[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel57[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel57[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel57[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel57[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel57[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel57[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel57[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel57[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel57[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel57[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel57[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel57[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel57[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel57[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel57[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel57[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel57[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel57[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel57[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel57[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel57),
		.Data_Out(add_k57_Data_Out),
		.Valid_Out(add_kernel57_Valid_Out)
	);
	Batch_Norm bn_kernel57(
		.Data_A(32'b00111110011110001000011101011100),
		.Data_B(32'b10111110110101001000100011000011),
		.Data_In(add_k57_Data_Out),
		.Valid_In(add_kernel57_Valid_Out),
		.Data_Out(bn57_Data_Out),
		.Valid_Out(bn57_Valid_Out)
	);
	Relu_Core rl_kernel57(
		.Data_In(bn57_Data_Out),
		.Valid_In(bn57_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*57-1:DATA_WIDHT*56]),
		.Valid_Out(rl57_Valid_Out)
	);
//////////KERNEL58//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111111011110111111101101100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110100000000101011110001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110111001010011110011000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111111001010000110011101000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111110000101011110111101101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111111000010110100100110001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111101110011101000000111101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111110101001110101110011011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110111100100110010011100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111110001001101000111001101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111110011011010101100100010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111111000000010001111001010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111101100111110000000001111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111110101000011000010110011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110000100110111100010100000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111101101111010101000010100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110101000110111001000001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111101111011011100000111011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111101001111010111010100101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111110011111001100000011000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110011110110000101010110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111111000011000001111000100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111110110011011001100111101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111110110110011111010011110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111110111101001111111100110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111011010001000001110111001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110101001010000010101111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111110101011101011001000001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111110011101100111000111100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110011000001011001110100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111110010111001111011000011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel58_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel58 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111110011001110100000101111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel58[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel58_Valid_Out)
	);
	Adder_32input add_k58(
		.Data1(Data_Out_Kernel58[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel58[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel58[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel58[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel58[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel58[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel58[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel58[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel58[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel58[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel58[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel58[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel58[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel58[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel58[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel58[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel58[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel58[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel58[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel58[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel58[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel58[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel58[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel58[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel58[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel58[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel58[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel58[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel58[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel58[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel58[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel58[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel58),
		.Data_Out(add_k58_Data_Out),
		.Valid_Out(add_kernel58_Valid_Out)
	);
	Batch_Norm bn_kernel58(
		.Data_A(32'b00111110011100100001111001101100),
		.Data_B(32'b10111110101100101001110001101111),
		.Data_In(add_k58_Data_Out),
		.Valid_In(add_kernel58_Valid_Out),
		.Data_Out(bn58_Data_Out),
		.Valid_Out(bn58_Valid_Out)
	);
	Relu_Core rl_kernel58(
		.Data_In(bn58_Data_Out),
		.Valid_In(bn58_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*58-1:DATA_WIDHT*57]),
		.Valid_Out(rl58_Valid_Out)
	);
//////////KERNEL59//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111110000101000001000100110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b10111110000001100001011111110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110101110000010001010011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110000111000010111000100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111110001011011001001001011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b00111110110010010000000101100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111101000111100011111100100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111110111101011110100000100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111111000111100111011001010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110011111001100011111110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111100110001101111100110101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111111000001010010011100110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111101100111000110110001001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111111010000100100100001010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111101100111010100000010000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111111000111000111010111111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111110000110100000101100001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111110001111101101010011111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111101010101100000101110100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111110110110010011011111000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111110110011010110000111101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111110100110001010100101100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111110110001100010101110100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111110100000111000010100000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111110000010011010001000010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111110001100001111111110101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111111000000011110001101000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111100111100101000011011110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111111001011100110000011010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111110011010110111111011001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111110100100011101000010100101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel59_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel59 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111110101000100010110101010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel59[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel59_Valid_Out)
	);
	Adder_32input add_k59(
		.Data1(Data_Out_Kernel59[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel59[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel59[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel59[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel59[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel59[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel59[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel59[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel59[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel59[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel59[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel59[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel59[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel59[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel59[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel59[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel59[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel59[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel59[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel59[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel59[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel59[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel59[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel59[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel59[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel59[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel59[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel59[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel59[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel59[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel59[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel59[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel59),
		.Data_Out(add_k59_Data_Out),
		.Valid_Out(add_kernel59_Valid_Out)
	);
	Batch_Norm bn_kernel59(
		.Data_A(32'b00111110010111011101011111011011),
		.Data_B(32'b00111110100011011111000001101001),
		.Data_In(add_k59_Data_Out),
		.Valid_In(add_kernel59_Valid_Out),
		.Data_Out(bn59_Data_Out),
		.Valid_Out(bn59_Valid_Out)
	);
	Relu_Core rl_kernel59(
		.Data_In(bn59_Data_Out),
		.Valid_In(bn59_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*59-1:DATA_WIDHT*58]),
		.Valid_Out(rl59_Valid_Out)
	);
//////////KERNEL60//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111111000101110010110010010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111101100110100000101001111111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110000100000011001010001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111111010001111100100100001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b10111110010000111110100001111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110001010010101110000011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111101110010111001101011011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111110100101111100111100101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110110001001110111110010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111110100001110010000111110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111110101011100110111100101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111101110110101111010010110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b00111110001101010010110010001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111110111010000011111001001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111111001011101101101001010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111100110010011110010100111110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111110101000011011111000001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110001001011011001100001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111111000001101101100100000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111111000011101100010001011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111101100000101110111000101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111101000010001100001010110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110000101010100100100111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111111001001110100001100110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111101010110101001010010110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110010000010100110011100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111101000111101000111110100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111100100000101001011111110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111110110000111010101000110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111111001000011101111110100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111110010000101010001011101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel60_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel60 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111110101101110110110110100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel60[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel60_Valid_Out)
	);
	Adder_32input add_k60(
		.Data1(Data_Out_Kernel60[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel60[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel60[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel60[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel60[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel60[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel60[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel60[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel60[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel60[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel60[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel60[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel60[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel60[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel60[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel60[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel60[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel60[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel60[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel60[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel60[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel60[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel60[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel60[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel60[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel60[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel60[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel60[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel60[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel60[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel60[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel60[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel60),
		.Data_Out(add_k60_Data_Out),
		.Valid_Out(add_kernel60_Valid_Out)
	);
	Batch_Norm bn_kernel60(
		.Data_A(32'b00111110011011111110000110101011),
		.Data_B(32'b10111111010100101000001111111000),
		.Data_In(add_k60_Data_Out),
		.Valid_In(add_kernel60_Valid_Out),
		.Data_Out(bn60_Data_Out),
		.Valid_Out(bn60_Valid_Out)
	);
	Relu_Core rl_kernel60(
		.Data_In(bn60_Data_Out),
		.Valid_In(bn60_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*60-1:DATA_WIDHT*59]),
		.Valid_Out(rl60_Valid_Out)
	);
//////////KERNEL61//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111101000010101001010011000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111110110100111011100100000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111111000000001011111111000000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111110100101001110011110110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111101101010111011001110110110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110100100100111111011000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111111000001000110010111011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111110101001011111000100010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110000111011011100101010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111110001110001110100101010100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111110100011011101101100101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111101101001110010000001011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111111000001011101110101000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111101111001010010101010000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111110100000010100111001011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111111000000000101110010001110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111100110100110001010111111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111110100111111100100011101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111110110001101100110010111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111101101101000100001110001100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b10111101101000010100111010011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111111010010001110111100011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111101101111100011110111100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b00111110110010110010000010000010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111101000001001101111000010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111110100100110101100100010101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111111000010100001000001110000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b10111110011110101011111010110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111111011110101100100011001000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111110110110010010001010010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111110010111000011100000010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel61_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel61 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111101110110101111110010101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel61[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel61_Valid_Out)
	);
	Adder_32input add_k61(
		.Data1(Data_Out_Kernel61[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel61[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel61[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel61[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel61[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel61[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel61[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel61[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel61[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel61[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel61[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel61[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel61[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel61[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel61[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel61[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel61[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel61[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel61[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel61[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel61[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel61[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel61[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel61[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel61[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel61[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel61[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel61[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel61[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel61[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel61[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel61[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel61),
		.Data_Out(add_k61_Data_Out),
		.Valid_Out(add_kernel61_Valid_Out)
	);
	Batch_Norm bn_kernel61(
		.Data_A(32'b00111110011001101011110010110001),
		.Data_B(32'b00111111100111010001001101110100),
		.Data_In(add_k61_Data_Out),
		.Valid_In(add_kernel61_Valid_Out),
		.Data_Out(bn61_Data_Out),
		.Valid_Out(bn61_Valid_Out)
	);
	Relu_Core rl_kernel61(
		.Data_In(bn61_Data_Out),
		.Valid_In(bn61_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*61-1:DATA_WIDHT*60]),
		.Valid_Out(rl61_Valid_Out)
	);
//////////KERNEL62//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110100100000101110101110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111110011000100011010000100111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111111000110100001010000101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b10111110001110001000000101010111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111110100010001011101010101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110101110001110101011001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111110011101001100111001011011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111111010101100101100001111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111110100000110000101010111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111111001011011110010100000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111101001101111101000100010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110011100000100100111010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110100110110011011111101001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111101000100010100011010101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b00111101110100011101101110010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111101001000101100001110101111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b10111111001011001001110110000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111111001011111000001100111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111110101011111000011000000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111110101010101010111101001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111101110100011111111101111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111110001000010110111111111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111110000001000111010111110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111110000001000000001000001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111101100110110000001010111101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b00111101001011111000111110000110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111110100001110000000111110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111110101101001111101101110010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111110001000000101010011111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b10111110101001011111001010001101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111111001100011010000111011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel62_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel62 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111111001010101010010100011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel62[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel62_Valid_Out)
	);
	Adder_32input add_k62(
		.Data1(Data_Out_Kernel62[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel62[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel62[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel62[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel62[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel62[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel62[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel62[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel62[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel62[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel62[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel62[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel62[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel62[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel62[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel62[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel62[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel62[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel62[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel62[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel62[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel62[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel62[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel62[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel62[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel62[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel62[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel62[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel62[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel62[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel62[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel62[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel62),
		.Data_Out(add_k62_Data_Out),
		.Valid_Out(add_kernel62_Valid_Out)
	);
	Batch_Norm bn_kernel62(
		.Data_A(32'b00111110011000000000110011011011),
		.Data_B(32'b10111110001011001110111111101100),
		.Data_In(add_k62_Data_Out),
		.Valid_In(add_kernel62_Valid_Out),
		.Data_Out(bn62_Data_Out),
		.Valid_Out(bn62_Valid_Out)
	);
	Relu_Core rl_kernel62(
		.Data_In(bn62_Data_Out),
		.Valid_In(bn62_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*62-1:DATA_WIDHT*61]),
		.Valid_Out(rl62_Valid_Out)
	);
//////////KERNEL63//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b10111110001100100011010000011110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111110100101100100001101111100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b00111110110000010001110111100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111101001000110000111000101011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111110110101011111010110111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110010100101111110110000100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b10111111000111110101001101000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b10111100101100010110000101010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b10111110000010010110111100111011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b00111101010101001011011110011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111101010111111110001101011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b00111110110010100011010000010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110010001001101110000111000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b10111110100101111100101100011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111111010011110101110101101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b10111110010001111001010011000101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111100100111011110011111000011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b00111111011111100111000011110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b10111110100001101100011110111001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b10111110010111111001011001010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111100110101001101110110100010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b00111110100001000101110010101010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b10111110100100001010111011101100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111110110111100101011001001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b00111111001111001010100010010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111010111011101100011001101110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b10111110111000110101011100010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111110100101000110101110010000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b00111110110111001111000010001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111110110111101110100000011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b00111101011011011000010000110101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel63_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel63 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111110000111111001111111100011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel63[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel63_Valid_Out)
	);
	Adder_32input add_k63(
		.Data1(Data_Out_Kernel63[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel63[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel63[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel63[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel63[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel63[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel63[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel63[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel63[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel63[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel63[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel63[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel63[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel63[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel63[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel63[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel63[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel63[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel63[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel63[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel63[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel63[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel63[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel63[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel63[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel63[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel63[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel63[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel63[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel63[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel63[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel63[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel63),
		.Data_Out(add_k63_Data_Out),
		.Valid_Out(add_kernel63_Valid_Out)
	);
	Batch_Norm bn_kernel63(
		.Data_A(32'b00111110100011010100110101110111),
		.Data_B(32'b00111111010110011101111110111101),
		.Data_In(add_k63_Data_Out),
		.Valid_In(add_kernel63_Valid_Out),
		.Data_Out(bn63_Data_Out),
		.Valid_Out(bn63_Valid_Out)
	);
	Relu_Core rl_kernel63(
		.Data_In(bn63_Data_Out),
		.Valid_In(bn63_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*63-1:DATA_WIDHT*62]),
		.Valid_Out(rl63_Valid_Out)
	);
//////////KERNEL64//////////
	Convolution2D_1x1_stride_1x1 CHANNEL1_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT-1:0]),
		.Kernel(32'b00111101100011010011110110001011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT-1:0]),
		.Valid_Out(channel1_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL2_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Kernel(32'b00111100011011010100111101101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*2-1:DATA_WIDHT*1]),
		.Valid_Out(channel2_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL3_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Kernel(32'b10111111000111101011101000011000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Valid_Out(channel3_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL4_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Kernel(32'b00111111000100101001011101101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Valid_Out(channel4_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL5_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Kernel(32'b00111110111100001001011011001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Valid_Out(channel5_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL6_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Kernel(32'b10111110110011010001100001110001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Valid_Out(channel6_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL7_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Kernel(32'b00111111001111011110101101010011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Valid_Out(channel7_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL8_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Kernel(32'b00111110101000100111100101010010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Valid_Out(channel8_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL9_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Kernel(32'b00111101101111011111000101000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Valid_Out(channel9_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL10_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Kernel(32'b10111110010011111010001101100001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Valid_Out(channel10_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL11_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Kernel(32'b10111101100001111111110100011010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Valid_Out(channel11_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL12_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Kernel(32'b10111111001110110000101101011111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Valid_Out(channel12_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL13_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Kernel(32'b10111110111000001101110001101101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Valid_Out(channel13_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL14_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Kernel(32'b00111101100000000110010000101000),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Valid_Out(channel14_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL15_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Kernel(32'b10111011001101101110010010001001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Valid_Out(channel15_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL16_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Kernel(32'b00111110000101010101111001001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Valid_Out(channel16_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL17_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Kernel(32'b00111101100000000111100101000001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Valid_Out(channel17_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL18_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Kernel(32'b10111110010111001111101011000111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Valid_Out(channel18_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL19_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Kernel(32'b00111110111111101011111011110100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Valid_Out(channel19_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL20_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Kernel(32'b00111111001001010100001000001111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Valid_Out(channel20_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL21_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Kernel(32'b00111110110010010001100001010110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Valid_Out(channel21_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL22_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Kernel(32'b10111110111000001101100111010001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Valid_Out(channel22_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL23_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Kernel(32'b00111110111111110111000111011100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Valid_Out(channel23_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL24_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Kernel(32'b10111101110010100001111000001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Valid_Out(channel24_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL25_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Kernel(32'b10111101100010001111101111011001),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Valid_Out(channel25_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL26_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Kernel(32'b10111111001000100001001110111010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Valid_Out(channel26_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL27_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Kernel(32'b00111110111111010010100001001010),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Valid_Out(channel27_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL28_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Kernel(32'b00111110101100000110001000110111),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Valid_Out(channel28_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL29_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Kernel(32'b10111101011001111100100011011101),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Valid_Out(channel29_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL30_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Kernel(32'b00111101110010001000010101100110),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Valid_Out(channel30_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL31_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Kernel(32'b10111101011011100000110010100100),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Valid_Out(channel31_Kernel64_Valid_Out)
	);
	Convolution2D_1x1_stride_1x1 CHANNEL32_Kernel64 (
		.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Kernel(32'b10111011101110000011010010110011),
		.Valid_In(Valid_In),
		.clk(clk),
		.rst(rst),
		.Data_Out(Data_Out_Kernel64[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_Out(channel32_Kernel64_Valid_Out)
	);
	Adder_32input add_k64(
		.Data1(Data_Out_Kernel64[DATA_WIDHT-1:0]),
		.Data2(Data_Out_Kernel64[DATA_WIDHT*2-1:DATA_WIDHT]),
		.Data3(Data_Out_Kernel64[DATA_WIDHT*3-1:DATA_WIDHT*2]),
		.Data4(Data_Out_Kernel64[DATA_WIDHT*4-1:DATA_WIDHT*3]),
		.Data5(Data_Out_Kernel64[DATA_WIDHT*5-1:DATA_WIDHT*4]),
		.Data6(Data_Out_Kernel64[DATA_WIDHT*6-1:DATA_WIDHT*5]),
		.Data7(Data_Out_Kernel64[DATA_WIDHT*7-1:DATA_WIDHT*6]),
		.Data8(Data_Out_Kernel64[DATA_WIDHT*8-1:DATA_WIDHT*7]),
		.Data9(Data_Out_Kernel64[DATA_WIDHT*9-1:DATA_WIDHT*8]),
		.Data10(Data_Out_Kernel64[DATA_WIDHT*10-1:DATA_WIDHT*9]),
		.Data11(Data_Out_Kernel64[DATA_WIDHT*11-1:DATA_WIDHT*10]),
		.Data12(Data_Out_Kernel64[DATA_WIDHT*12-1:DATA_WIDHT*11]),
		.Data13(Data_Out_Kernel64[DATA_WIDHT*13-1:DATA_WIDHT*12]),
		.Data14(Data_Out_Kernel64[DATA_WIDHT*14-1:DATA_WIDHT*13]),
		.Data15(Data_Out_Kernel64[DATA_WIDHT*15-1:DATA_WIDHT*14]),
		.Data16(Data_Out_Kernel64[DATA_WIDHT*16-1:DATA_WIDHT*15]),
		.Data17(Data_Out_Kernel64[DATA_WIDHT*17-1:DATA_WIDHT*16]),
		.Data18(Data_Out_Kernel64[DATA_WIDHT*18-1:DATA_WIDHT*17]),
		.Data19(Data_Out_Kernel64[DATA_WIDHT*19-1:DATA_WIDHT*18]),
		.Data20(Data_Out_Kernel64[DATA_WIDHT*20-1:DATA_WIDHT*19]),
		.Data21(Data_Out_Kernel64[DATA_WIDHT*21-1:DATA_WIDHT*20]),
		.Data22(Data_Out_Kernel64[DATA_WIDHT*22-1:DATA_WIDHT*21]),
		.Data23(Data_Out_Kernel64[DATA_WIDHT*23-1:DATA_WIDHT*22]),
		.Data24(Data_Out_Kernel64[DATA_WIDHT*24-1:DATA_WIDHT*23]),
		.Data25(Data_Out_Kernel64[DATA_WIDHT*25-1:DATA_WIDHT*24]),
		.Data26(Data_Out_Kernel64[DATA_WIDHT*26-1:DATA_WIDHT*25]),
		.Data27(Data_Out_Kernel64[DATA_WIDHT*27-1:DATA_WIDHT*26]),
		.Data28(Data_Out_Kernel64[DATA_WIDHT*28-1:DATA_WIDHT*27]),
		.Data29(Data_Out_Kernel64[DATA_WIDHT*29-1:DATA_WIDHT*28]),
		.Data30(Data_Out_Kernel64[DATA_WIDHT*30-1:DATA_WIDHT*29]),
		.Data31(Data_Out_Kernel64[DATA_WIDHT*31-1:DATA_WIDHT*30]),
		.Data32(Data_Out_Kernel64[DATA_WIDHT*32-1:DATA_WIDHT*31]),
		.Valid_In(add_kernel64),
		.Data_Out(add_k64_Data_Out),
		.Valid_Out(add_kernel64_Valid_Out)
	);
	Batch_Norm bn_kernel64(
		.Data_A(32'b00111110011101011011101000111011),
		.Data_B(32'b00111111100001101101000010101110),
		.Data_In(add_k64_Data_Out),
		.Valid_In(add_kernel64_Valid_Out),
		.Data_Out(bn64_Data_Out),
		.Valid_Out(bn64_Valid_Out)
	);
	Relu_Core rl_kernel64(
		.Data_In(bn64_Data_Out),
		.Valid_In(bn64_Valid_Out),
		.Data_Out(Data_Out[DATA_WIDHT*64-1:DATA_WIDHT*63]),
		.Valid_Out(rl64_Valid_Out)
	);

endmodule