module Depthwise_Part1_Separable_32CHANNEL_Layer4 #(
    parameter DATA_WIDHT = 32, 
    parameter IMG_WIDHT = 44,
    parameter IMG_HEIGHT =44
)
(
    input [DATA_WIDHT*32-1:0] Data_In,
    input clk,
    input rst,
    input Valid_In,
    output [DATA_WIDHT*32-1:0] Data_Out,
    output Valid_Out

);
    wire CHANNEL1_Valid_Out, CHANNEL2_Valid_Out, CHANNEL3_Valid_Out, CHANNEL4_Valid_Out, CHANNEL5_Valid_Out, CHANNEL6_Valid_Out, CHANNEL7_Valid_Out, CHANNEL8_Valid_Out, CHANNEL9_Valid_Out, CHANNEL10_Valid_Out, CHANNEL11_Valid_Out, CHANNEL12_Valid_Out, CHANNEL13_Valid_Out, CHANNEL14_Valid_Out, CHANNEL15_Valid_Out, CHANNEL16_Valid_Out, CHANNEL17_Valid_Out, CHANNEL18_Valid_Out, CHANNEL19_Valid_Out, CHANNEL20_Valid_Out, CHANNEL21_Valid_Out, CHANNEL22_Valid_Out, CHANNEL23_Valid_Out, CHANNEL24_Valid_Out,CHANNEL25_Valid_Out,CHANNEL26_Valid_Out,CHANNEL27_Valid_Out,CHANNEL28_Valid_Out,CHANNEL29_Valid_Out,CHANNEL30_Valid_Out,CHANNEL31_Valid_Out,CHANNEL32_Valid_Out;

	assign Valid_Out= CHANNEL1_Valid_Out & CHANNEL2_Valid_Out & CHANNEL3_Valid_Out & CHANNEL4_Valid_Out & CHANNEL5_Valid_Out & CHANNEL6_Valid_Out & CHANNEL7_Valid_Out & CHANNEL8_Valid_Out & CHANNEL9_Valid_Out & CHANNEL10_Valid_Out & CHANNEL11_Valid_Out & CHANNEL12_Valid_Out & CHANNEL13_Valid_Out & CHANNEL14_Valid_Out & CHANNEL15_Valid_Out & CHANNEL16_Valid_Out & CHANNEL17_Valid_Out & CHANNEL18_Valid_Out & CHANNEL19_Valid_Out & CHANNEL20_Valid_Out & CHANNEL21_Valid_Out & CHANNEL22_Valid_Out& CHANNEL23_Valid_Out& CHANNEL24_Valid_Out&CHANNEL25_Valid_Out&CHANNEL26_Valid_Out&CHANNEL27_Valid_Out&CHANNEL28_Valid_Out&CHANNEL29_Valid_Out&CHANNEL30_Valid_Out&CHANNEL31_Valid_Out&CHANNEL32_Valid_Out;
		Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL1 (
			.Data_In(Data_In[DATA_WIDHT-1:0]),
			.Kernel0(32'b10111110000011011101011110101000),
			.Kernel1(32'b00111111000000001111110100000001),
			.Kernel2(32'b00111110100100110111000100111101),
			.Kernel3(32'b00111110001101011110000101101011),
			.Kernel4(32'b10111110011110000010011100111011),
			.Kernel5(32'b00111101101100101010000001011011),
			.Kernel6(32'b10111111000010001101000011101110),
			.Kernel7(32'b10111111010101100011010001010000),
			.Kernel8(32'b10111111000001100000110110101111),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT-1:0]),
			.Valid_Out(CHANNEL1_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL2 (
			.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
			.Kernel0(32'b10111110101101000001111101110010),
			.Kernel1(32'b10111110110011010101001010110011),
			.Kernel2(32'b10111110110001111001111111011001),
			.Kernel3(32'b10111110110001101101000001000000),
			.Kernel4(32'b10111101111101010001010001001001),
			.Kernel5(32'b00111101011101011111001001010100),
			.Kernel6(32'b00111110111000011011100000100010),
			.Kernel7(32'b00111110111000001001010101101101),
			.Kernel8(32'b00111111000110101000001100001101),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*2-1:DATA_WIDHT]),
			.Valid_Out(CHANNEL2_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL3 (
			.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
			.Kernel0(32'b00111110111011110000000010010011),
			.Kernel1(32'b00111111001101100000100011111001),
			.Kernel2(32'b00111111000101000011111011111111),
			.Kernel3(32'b10111100111010001101111011100001),
			.Kernel4(32'b10111101110101010101010010000001),
			.Kernel5(32'b10111110100110001010001100001100),
			.Kernel6(32'b10111111001111100111000011100011),
			.Kernel7(32'b10111110011010011110010110010110),
			.Kernel8(32'b10111111000111001100011001001001),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*3-1:DATA_WIDHT*2]),
			.Valid_Out(CHANNEL3_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL4 (
			.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
			.Kernel0(32'b00111110111011100001100011100111),
			.Kernel1(32'b10111110110101001101110000100001),
			.Kernel2(32'b00111111011001001001100111100010),
			.Kernel3(32'b00111101111011111100010010101001),
			.Kernel4(32'b10111110111110111100001111001110),
			.Kernel5(32'b00111100001110011100001011011100),
			.Kernel6(32'b10111110100100000111101101001000),
			.Kernel7(32'b10111111000000011101001111011111),
			.Kernel8(32'b10111101110000011000101100001011),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*4-1:DATA_WIDHT*3]),
			.Valid_Out(CHANNEL4_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL5 (
			.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
			.Kernel0(32'b00111111010111011111011011001010),
			.Kernel1(32'b00111110001101101001010011100101),
			.Kernel2(32'b00111111000010110011000010001010),
			.Kernel3(32'b10111110100110000001100010101010),
			.Kernel4(32'b00111110100010101100011101111101),
			.Kernel5(32'b10111100001000001001101110001011),
			.Kernel6(32'b10111010000111010111001001100100),
			.Kernel7(32'b00111111000001100001101100101000),
			.Kernel8(32'b00111110000000111111001010100001),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*5-1:DATA_WIDHT*4]),
			.Valid_Out(CHANNEL5_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL6 (
			.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
			.Kernel0(32'b00111111000001100000001100011010),
			.Kernel1(32'b00111111001010011110000010100000),
			.Kernel2(32'b00111111010010110001111000100000),
			.Kernel3(32'b00111101010010010001100101010111),
			.Kernel4(32'b10111101111000010000001000110011),
			.Kernel5(32'b10111101110011000011110100001101),
			.Kernel6(32'b10111110001111100001011000011101),
			.Kernel7(32'b00111110001001101001011110101010),
			.Kernel8(32'b10111110111010101011100001010010),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*6-1:DATA_WIDHT*5]),
			.Valid_Out(CHANNEL6_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL7 (
			.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
			.Kernel0(32'b10111101111010000101000100101000),
			.Kernel1(32'b00111110001110111001111000000110),
			.Kernel2(32'b10111110100111010110110011001101),
			.Kernel3(32'b00111110000011001000110011100100),
			.Kernel4(32'b00111100001001110100101110110111),
			.Kernel5(32'b00111111000110010100011000001001),
			.Kernel6(32'b00111110101110001011000110010001),
			.Kernel7(32'b00111111000100100100001000001100),
			.Kernel8(32'b00111111000001000100001000011010),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*7-1:DATA_WIDHT*6]),
			.Valid_Out(CHANNEL7_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL8 (
			.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
			.Kernel0(32'b00111110111011000011001011010001),
			.Kernel1(32'b10111110010000111011101010010111),
			.Kernel2(32'b00111110111010011010101110101010),
			.Kernel3(32'b00111111001000100111111010110100),
			.Kernel4(32'b00111101001010110000011100000100),
			.Kernel5(32'b00111110111110100000100010110010),
			.Kernel6(32'b00111110111100100101010000001010),
			.Kernel7(32'b10111110000101111111011100010111),
			.Kernel8(32'b00111110100000111110100011110111),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*8-1:DATA_WIDHT*7]),
			.Valid_Out(CHANNEL8_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL9 (
			.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
			.Kernel0(32'b00111101100010011010111110000000),
			.Kernel1(32'b10111110111010100010101110011111),
			.Kernel2(32'b10111110110001111111110101111000),
			.Kernel3(32'b00111110111001011001100010010111),
			.Kernel4(32'b00111110100000111101110000111111),
			.Kernel5(32'b00111110110000111110010100111110),
			.Kernel6(32'b00111110010000110000110110001100),
			.Kernel7(32'b00111110001010111111010000110000),
			.Kernel8(32'b00111111001101100100110010111100),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*9-1:DATA_WIDHT*8]),
			.Valid_Out(CHANNEL9_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL10 (
			.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
			.Kernel0(32'b00111111001010011011011101111010),
			.Kernel1(32'b00111110001011000011001110010000),
			.Kernel2(32'b00111110100000110100101100001101),
			.Kernel3(32'b00111111000010001111100000100111),
			.Kernel4(32'b00111100111010001011100100011100),
			.Kernel5(32'b10111110010111000111010010111100),
			.Kernel6(32'b10111110000101111111110010110110),
			.Kernel7(32'b00111110111011001011000000011010),
			.Kernel8(32'b10111110011000100111101000000110),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*10-1:DATA_WIDHT*9]),
			.Valid_Out(CHANNEL10_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL11 (
			.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
			.Kernel0(32'b10111110111110010001110101101011),
			.Kernel1(32'b10111111000001001010001101101111),
			.Kernel2(32'b10111111000100110010101011101010),
			.Kernel3(32'b00111110110111001100111101111001),
			.Kernel4(32'b00111110111010110001111010000111),
			.Kernel5(32'b00111110011001001001011101111011),
			.Kernel6(32'b00111110101000010011000111111000),
			.Kernel7(32'b00111111000111110111011010110101),
			.Kernel8(32'b00111110000011111000111010110111),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*11-1:DATA_WIDHT*10]),
			.Valid_Out(CHANNEL11_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL12 (
			.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
			.Kernel0(32'b00111101111101110111111001111001),
			.Kernel1(32'b00111111000011100111110000010110),
			.Kernel2(32'b00111100000101110111000011000011),
			.Kernel3(32'b10111110000101010110000011000100),
			.Kernel4(32'b10111110100010111111011001110101),
			.Kernel5(32'b00111110100001010010000001110111),
			.Kernel6(32'b00111111000111011011011101011100),
			.Kernel7(32'b00111111001001110001000001101111),
			.Kernel8(32'b00111110100100100001000001000111),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*12-1:DATA_WIDHT*11]),
			.Valid_Out(CHANNEL12_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL13 (
			.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
			.Kernel0(32'b00111110000011101011010011001000),
			.Kernel1(32'b10111110100110111101110100101111),
			.Kernel2(32'b10111110010101010011010010110110),
			.Kernel3(32'b00111111001100011011011011110010),
			.Kernel4(32'b10111100011010011010011010111110),
			.Kernel5(32'b10111101000000111111011100011000),
			.Kernel6(32'b00111101111000011110010011110101),
			.Kernel7(32'b10111111000101000101010111010100),
			.Kernel8(32'b10111110111010111011101010101111),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*13-1:DATA_WIDHT*12]),
			.Valid_Out(CHANNEL13_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL14 (
			.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
			.Kernel0(32'b10111111010011111000111000111111),
			.Kernel1(32'b10111110110011010111110011000101),
			.Kernel2(32'b10111111011000000001000001011110),
			.Kernel3(32'b10111111000000001110101001011110),
			.Kernel4(32'b10111110001111001110111011101010),
			.Kernel5(32'b10111110110010110001110100111110),
			.Kernel6(32'b00111110011001011010101010011101),
			.Kernel7(32'b00111110101011010000100000100100),
			.Kernel8(32'b10111110110011010101011011111110),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*14-1:DATA_WIDHT*13]),
			.Valid_Out(CHANNEL14_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL15 (
			.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
			.Kernel0(32'b00111110111001111001110111011011),
			.Kernel1(32'b00111110110000100101100111010010),
			.Kernel2(32'b00111111000001000111011111111101),
			.Kernel3(32'b00111110011000110110001001111011),
			.Kernel4(32'b10111110111011011011011000011000),
			.Kernel5(32'b10111111000110001001110100001111),
			.Kernel6(32'b10111101001011101010010001101111),
			.Kernel7(32'b10111110101010000111110001100000),
			.Kernel8(32'b00111101101111100101110010110110),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*15-1:DATA_WIDHT*14]),
			.Valid_Out(CHANNEL15_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL16 (
			.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
			.Kernel0(32'b00111110001000001101000111010011),
			.Kernel1(32'b00111110000100000011011111101100),
			.Kernel2(32'b00111110101010100011100000010111),
			.Kernel3(32'b00111111000110000011011000001010),
			.Kernel4(32'b00111110110100000011110101000000),
			.Kernel5(32'b00111110111010101010110110010001),
			.Kernel6(32'b00111110100000101101101100110101),
			.Kernel7(32'b10111110011101000000111111000011),
			.Kernel8(32'b00111101000001110001000010001001),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*16-1:DATA_WIDHT*15]),
			.Valid_Out(CHANNEL16_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL17 (
			.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
			.Kernel0(32'b10111101100001111001011111100000),
			.Kernel1(32'b10111110101001000000010110011001),
			.Kernel2(32'b00111110000001000111000101011111),
			.Kernel3(32'b00111101010011111110111011010100),
			.Kernel4(32'b00111100101010111011001010101110),
			.Kernel5(32'b00111101110111111100010100010111),
			.Kernel6(32'b00111111001110001100000100001001),
			.Kernel7(32'b00111111000000000011000101100001),
			.Kernel8(32'b00111110111111111011011101110010),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*17-1:DATA_WIDHT*16]),
			.Valid_Out(CHANNEL17_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL18 (
			.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
			.Kernel0(32'b10111101000101010100111101111110),
			.Kernel1(32'b00111011001001110010011101100100),
			.Kernel2(32'b10111111000010100111000001011110),
			.Kernel3(32'b00111111000110001000011101100010),
			.Kernel4(32'b00111111010101010011001000001110),
			.Kernel5(32'b00111100011110000101101011010011),
			.Kernel6(32'b00111100110101011000010111010111),
			.Kernel7(32'b10111110001101010001010010100101),
			.Kernel8(32'b10111110110100000010101000101110),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*18-1:DATA_WIDHT*17]),
			.Valid_Out(CHANNEL18_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL19 (
			.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
			.Kernel0(32'b00111110110000011011110000001001),
			.Kernel1(32'b00111111000001000001001000111101),
			.Kernel2(32'b10111101011101011001001011010101),
			.Kernel3(32'b10111101110101101000100001001001),
			.Kernel4(32'b10111110001101111011111001010110),
			.Kernel5(32'b10111101110101111001111000111111),
			.Kernel6(32'b10111110110001011010001001101101),
			.Kernel7(32'b10111110101101101010101111010101),
			.Kernel8(32'b10111111011011011001001100011101),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*19-1:DATA_WIDHT*18]),
			.Valid_Out(CHANNEL19_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL20 (
			.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
			.Kernel0(32'b10111110101101100101000111011111),
			.Kernel1(32'b10111101001010100100101111100011),
			.Kernel2(32'b10111101111100100001100000000001),
			.Kernel3(32'b10111111000000000011001011101101),
			.Kernel4(32'b10111110110000011100000000100010),
			.Kernel5(32'b10111110100001111111000001100111),
			.Kernel6(32'b00111110101100011110000100011101),
			.Kernel7(32'b00111111001010111011010011001001),
			.Kernel8(32'b00111110100110110100010110110110),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*20-1:DATA_WIDHT*19]),
			.Valid_Out(CHANNEL20_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL21 (
			.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
			.Kernel0(32'b00111111000100011101000110010000),
			.Kernel1(32'b00111110010100000000110000100010),
			.Kernel2(32'b00111111000111111000010111100100),
			.Kernel3(32'b10111110010100110010010110111011),
			.Kernel4(32'b00111110111001010111111011011010),
			.Kernel5(32'b00111110111011010000011111001100),
			.Kernel6(32'b00111101010101110000010101110111),
			.Kernel7(32'b10111110010011010101000010011100),
			.Kernel8(32'b10111100111100101111101101111010),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*21-1:DATA_WIDHT*20]),
			.Valid_Out(CHANNEL21_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL22 (
			.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
			.Kernel0(32'b10111011101011111100100001111010),
			.Kernel1(32'b00111101001001011100110111110001),
			.Kernel2(32'b00111101100001110110101011011110),
			.Kernel3(32'b10111111000101011010111010010001),
			.Kernel4(32'b10111110101111101101100100111000),
			.Kernel5(32'b10111110111011010100011110011101),
			.Kernel6(32'b10111110001111011001000011100000),
			.Kernel7(32'b10111110010100110001000111101000),
			.Kernel8(32'b10111111001011001100001101110001),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*22-1:DATA_WIDHT*21]),
			.Valid_Out(CHANNEL22_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL23 (
			.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
			.Kernel0(32'b00111110110110101001010000001100),
			.Kernel1(32'b00111110001110001011100110000000),
			.Kernel2(32'b00111111001000001011001100111101),
			.Kernel3(32'b10111110100111100011010101111101),
			.Kernel4(32'b10111110111000110001011000110101),
			.Kernel5(32'b00111101111011001001110110110010),
			.Kernel6(32'b00111110110100100110110000101001),
			.Kernel7(32'b00111110001100010111111110001011),
			.Kernel8(32'b00111110111100000011011000100100),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*23-1:DATA_WIDHT*22]),
			.Valid_Out(CHANNEL23_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL24 (
			.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
			.Kernel0(32'b10111111001011000101011111110110),
			.Kernel1(32'b10111110011010110000010010000110),
			.Kernel2(32'b10111111011011010011101011100111),
			.Kernel3(32'b00111110000110010111010010011011),
			.Kernel4(32'b00111110000101101011010100110001),
			.Kernel5(32'b10111110001110000001100101101111),
			.Kernel6(32'b00111110100001101101100001101110),
			.Kernel7(32'b00111111000000110111111010000111),
			.Kernel8(32'b00111110011111000000100001101010),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*24-1:DATA_WIDHT*23]),
			.Valid_Out(CHANNEL24_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL25 (
			.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
			.Kernel0(32'b00111110101101111001111010100010),
			.Kernel1(32'b00111111000001001100001000111110),
			.Kernel2(32'b00111111000110100010011111001010),
			.Kernel3(32'b10111111001110111100111111010100),
			.Kernel4(32'b10111110010010011101000011000100),
			.Kernel5(32'b10111111001001001011100110100101),
			.Kernel6(32'b10111101010100110010100011101110),
			.Kernel7(32'b00111110101100110001110000110111),
			.Kernel8(32'b10111101010000110111001010001010),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*25-1:DATA_WIDHT*24]),
			.Valid_Out(CHANNEL25_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL26 (
			.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
			.Kernel0(32'b10111110111101111010010001101111),
			.Kernel1(32'b00111110101010010110101001010010),
			.Kernel2(32'b10111110110110010000010010100000),
			.Kernel3(32'b10111110000010010110010011001010),
			.Kernel4(32'b00111100111100100011000000011110),
			.Kernel5(32'b10111110110000010000011000001000),
			.Kernel6(32'b00111100100010001101011100101110),
			.Kernel7(32'b00111111000011101111111000010001),
			.Kernel8(32'b00111110110000100111000001111011),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*26-1:DATA_WIDHT*25]),
			.Valid_Out(CHANNEL26_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL27 (
			.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
			.Kernel0(32'b10111110101100101100010000100000),
			.Kernel1(32'b10111111001100110101111000001011),
			.Kernel2(32'b10111101111111010110010001001111),
			.Kernel3(32'b10111110000101011100101011011010),
			.Kernel4(32'b00111110010011101100001011110101),
			.Kernel5(32'b10111110000001010100100100111110),
			.Kernel6(32'b10111111000010010000001110110011),
			.Kernel7(32'b10111101101000000010110100010001),
			.Kernel8(32'b10111110111010110000001110111010),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*27-1:DATA_WIDHT*26]),
			.Valid_Out(CHANNEL27_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL28 (
			.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
			.Kernel0(32'b00111111000001101101111000101110),
			.Kernel1(32'b00111110011001111100011110100010),
			.Kernel2(32'b10111101100011000010111111000001),
			.Kernel3(32'b00111110111100001111110001001111),
			.Kernel4(32'b00111111001111001101100001100101),
			.Kernel5(32'b00111110111010110001000111111001),
			.Kernel6(32'b00111110101001001101101100011110),
			.Kernel7(32'b00111110000110111010000100110010),
			.Kernel8(32'b10111110111101000000011010000011),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*28-1:DATA_WIDHT*27]),
			.Valid_Out(CHANNEL28_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL29 (
			.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
			.Kernel0(32'b10111111010110111111101001000010),
			.Kernel1(32'b10111110010111110001111110010011),
			.Kernel2(32'b10111111001110000111111110001000),
			.Kernel3(32'b00111011111001101110010010111000),
			.Kernel4(32'b00111110010110101010011000110100),
			.Kernel5(32'b00111101011100111110110110001011),
			.Kernel6(32'b10111101100101111111001011010110),
			.Kernel7(32'b10111101011011010011010011001011),
			.Kernel8(32'b10111101101110100000101011101111),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*29-1:DATA_WIDHT*28]),
			.Valid_Out(CHANNEL29_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL30 (
			.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
			.Kernel0(32'b10111101000010010001010101010010),
			.Kernel1(32'b00111011110100101101101100011001),
			.Kernel2(32'b00111101001110010111100011001010),
			.Kernel3(32'b00111101101011000010001011000100),
			.Kernel4(32'b00111111011000011001101000011100),
			.Kernel5(32'b00111110110111001101001100000000),
			.Kernel6(32'b00111101111010011001100001111100),
			.Kernel7(32'b00111110100001100111101111011110),
			.Kernel8(32'b00111101010110001010101101111101),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*30-1:DATA_WIDHT*29]),
			.Valid_Out(CHANNEL30_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL31 (
			.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
			.Kernel0(32'b00111111001101001101010010101001),
			.Kernel1(32'b00111111000010000100011101000000),
			.Kernel2(32'b00111110100100110010100100110110),
			.Kernel3(32'b00111110111110001010001000010101),
			.Kernel4(32'b00111110110101000011111010000101),
			.Kernel5(32'b00111110111100000011111000101110),
			.Kernel6(32'b00111110010110001101011111110011),
			.Kernel7(32'b10111110010100010111001011010000),
			.Kernel8(32'b10111101010100011001101010001011),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*31-1:DATA_WIDHT*30]),
			.Valid_Out(CHANNEL31_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL32 (
			.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
			.Kernel0(32'b10111101110100010011001010100011),
			.Kernel1(32'b00111111001000100000111011100101),
			.Kernel2(32'b00111110111011110011110000001110),
			.Kernel3(32'b10111110100100000100100110111101),
			.Kernel4(32'b10111101101010101100111101110111),
			.Kernel5(32'b00111101001000110100111010100000),
			.Kernel6(32'b00111001011001000011101010001001),
			.Kernel7(32'b10111111010011010011100000110110),
			.Kernel8(32'b10111110101110101011010011000111),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*32-1:DATA_WIDHT*31]),
			.Valid_Out(CHANNEL32_Valid_Out)
		);

    
endmodule