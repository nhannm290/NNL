module Depthwise_Part1_Separable_16CHANNEL_Layer4  #(
    parameter DATA_WIDHT = 32, 
    parameter IMG_WIDHT = 44,
    parameter IMG_HEIGHT =44
)
(
    input [DATA_WIDHT*16-1:0] Data_In,
    input clk,
    input rst,
    input Valid_In,
    output [DATA_WIDHT*16-1:0] Data_Out,
    output Valid_Out

);

    wire CHANNEL1_Valid_Out, CHANNEL2_Valid_Out, CHANNEL3_Valid_Out, CHANNEL4_Valid_Out, CHANNEL5_Valid_Out, CHANNEL6_Valid_Out, CHANNEL7_Valid_Out, CHANNEL8_Valid_Out, CHANNEL9_Valid_Out, CHANNEL10_Valid_Out, CHANNEL11_Valid_Out, CHANNEL12_Valid_Out, CHANNEL13_Valid_Out, CHANNEL14_Valid_Out, CHANNEL15_Valid_Out, CHANNEL16_Valid_Out;

	assign Valid_Out= CHANNEL1_Valid_Out & CHANNEL2_Valid_Out & CHANNEL3_Valid_Out & CHANNEL4_Valid_Out & CHANNEL5_Valid_Out & CHANNEL6_Valid_Out & CHANNEL7_Valid_Out & CHANNEL8_Valid_Out & CHANNEL9_Valid_Out & CHANNEL10_Valid_Out & CHANNEL11_Valid_Out & CHANNEL12_Valid_Out & CHANNEL13_Valid_Out & CHANNEL14_Valid_Out & CHANNEL15_Valid_Out & CHANNEL16_Valid_Out;


	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL1 (
			.Data_In(Data_In[DATA_WIDHT-1:0]),
			.Kernel0(32'b00111110001000110101100001101011),
			.Kernel1(32'b00111111000100101001011001000000),
			.Kernel2(32'b10111101011111001111010111000000),
			.Kernel3(32'b10111110011101100101101111101100),
			.Kernel4(32'b10111110100001101101010101010111),
			.Kernel5(32'b10111101001100011000101100100111),
			.Kernel6(32'b10111111011000101110011111111100),
			.Kernel7(32'b10111111001010011001001100001100),
			.Kernel8(32'b10111110011101010000000010010111),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT-1:0]),
			.Valid_Out(CHANNEL1_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL2 (
			.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
			.Kernel0(32'b00111111001010010101110011011101),
			.Kernel1(32'b00111101110100100011000110110001),
			.Kernel2(32'b00111110111011101010100011000110),
			.Kernel3(32'b00111101010000111000001001011000),
			.Kernel4(32'b10111111000110001110110011100010),
			.Kernel5(32'b00111110010010000010101110001001),
			.Kernel6(32'b00111110100110111100100011010001),
			.Kernel7(32'b10111111000011111110000000100010),
			.Kernel8(32'b00111110100101110110110100011110),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*2-1:DATA_WIDHT]),
			.Valid_Out(CHANNEL2_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL3 (
			.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
			.Kernel0(32'b00111101100100100011100101110001),
			.Kernel1(32'b10111101100001111100000110111001),
			.Kernel2(32'b00111110110110111010101000100110),
			.Kernel3(32'b10111110101111010011001010110011),
			.Kernel4(32'b00111110000101111111110000100011),
			.Kernel5(32'b10111111000100001111100010011110),
			.Kernel6(32'b10111110101110110010010100010010),
			.Kernel7(32'b10111111000000111101100100001111),
			.Kernel8(32'b10111110100111101011000000100001),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*3-1:DATA_WIDHT*2]),
			.Valid_Out(CHANNEL3_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL4 (
			.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
			.Kernel0(32'b10111111010011111101000100001011),
			.Kernel1(32'b10111111000111010010011000011100),
			.Kernel2(32'b10111110100010001101010011101001),
			.Kernel3(32'b00111110000001110110110011001110),
			.Kernel4(32'b00111111000010110111001001000101),
			.Kernel5(32'b10111110000111111000100011111001),
			.Kernel6(32'b00111110111010111001001000000101),
			.Kernel7(32'b00111110100100100001100100111100),
			.Kernel8(32'b00111110100101010111110101101000),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*4-1:DATA_WIDHT*3]),
			.Valid_Out(CHANNEL4_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL5 (
			.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
			.Kernel0(32'b00111110111111011101001001110010),
			.Kernel1(32'b00111110110111000001100001001000),
			.Kernel2(32'b00111110101011111000101011010110),
			.Kernel3(32'b00111110000000010110110111000011),
			.Kernel4(32'b10111110100110011000010110001010),
			.Kernel5(32'b00111110111101110011010011111010),
			.Kernel6(32'b00111100100101001011100110001100),
			.Kernel7(32'b00111110110111101000101000011010),
			.Kernel8(32'b00111110101010101010101101010101),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*5-1:DATA_WIDHT*4]),
			.Valid_Out(CHANNEL5_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL6 (
			.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
			.Kernel0(32'b10111110110101010110100011001010),
			.Kernel1(32'b10111110011101000110101010100110),
			.Kernel2(32'b10111110000010110101111011110011),
			.Kernel3(32'b10111110111000100000101010111010),
			.Kernel4(32'b10111110010110111111101100000111),
			.Kernel5(32'b10111101001001100101010100110110),
			.Kernel6(32'b10111110100011000100101010011100),
			.Kernel7(32'b10111101000100001101011001100010),
			.Kernel8(32'b10111100100101000011000100111010),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*6-1:DATA_WIDHT*5]),
			.Valid_Out(CHANNEL6_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL7 (
			.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
			.Kernel0(32'b10111110100010101011101101011100),
			.Kernel1(32'b00111110001110010011111010110010),
			.Kernel2(32'b00111101000010111010110101000000),
			.Kernel3(32'b10111101100100101000011111111011),
			.Kernel4(32'b00111110001010110100110100101000),
			.Kernel5(32'b10111100111111101110111101010010),
			.Kernel6(32'b10111111100011001110101101101101),
			.Kernel7(32'b10111111010110111111010001010110),
			.Kernel8(32'b10111111000111010010110010101110),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*7-1:DATA_WIDHT*6]),
			.Valid_Out(CHANNEL7_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL8 (
			.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
			.Kernel0(32'b10111101001100110110110100001000),
			.Kernel1(32'b00111110011010000110011001001010),
			.Kernel2(32'b10111110100001111111000010101110),
			.Kernel3(32'b10111110111111000010001010011010),
			.Kernel4(32'b10111110100000100101010100011011),
			.Kernel5(32'b10111110111110101011101100110000),
			.Kernel6(32'b00111110011001100010010000110100),
			.Kernel7(32'b00111110110010101010100001101000),
			.Kernel8(32'b10111110001101111011000011100110),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*8-1:DATA_WIDHT*7]),
			.Valid_Out(CHANNEL8_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL9 (
			.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
			.Kernel0(32'b10111110111011110011000000110100),
			.Kernel1(32'b00111101100101011010011001011010),
			.Kernel2(32'b10111110101110001101000001100110),
			.Kernel3(32'b10111110110101101000101101110001),
			.Kernel4(32'b00111101001100010000010001111011),
			.Kernel5(32'b10111111000000101110000101101001),
			.Kernel6(32'b10111110110010001010010001010111),
			.Kernel7(32'b10111110110000010111011101111110),
			.Kernel8(32'b10111110011100010000111000010111),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*9-1:DATA_WIDHT*8]),
			.Valid_Out(CHANNEL9_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL10 (
			.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
			.Kernel0(32'b10111110100000110001111111101001),
			.Kernel1(32'b10111110101010100111011011001100),
			.Kernel2(32'b00111011111101100110100101101000),
			.Kernel3(32'b10111111001101000001110111001110),
			.Kernel4(32'b10111110000111001110110010100101),
			.Kernel5(32'b10111110100000110110111001001100),
			.Kernel6(32'b10111111000010011110001011101110),
			.Kernel7(32'b00111100100101001101110011000101),
			.Kernel8(32'b10111110110101010000100000001101),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*10-1:DATA_WIDHT*9]),
			.Valid_Out(CHANNEL10_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL11 (
			.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
			.Kernel0(32'b00111111011110010001000100100100),
			.Kernel1(32'b00111100011000101100001111100000),
			.Kernel2(32'b00111111001111101100100010111111),
			.Kernel3(32'b00111110100101111010011001001110),
			.Kernel4(32'b10111110101000110001001000000000),
			.Kernel5(32'b00111110001010111001010000100101),
			.Kernel6(32'b10111101101100001110101011001010),
			.Kernel7(32'b10111110111101100011001011000010),
			.Kernel8(32'b00111110101100101100101011010100),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*11-1:DATA_WIDHT*10]),
			.Valid_Out(CHANNEL11_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL12 (
			.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
			.Kernel0(32'b10111110101010110101101110011010),
			.Kernel1(32'b00111110100001111110110001100001),
			.Kernel2(32'b10111110000000010001010110110101),
			.Kernel3(32'b10111110111011000110101111011000),
			.Kernel4(32'b00111100100011111101110001100000),
			.Kernel5(32'b10111111000000001011010101100111),
			.Kernel6(32'b10111110010010001010110000111110),
			.Kernel7(32'b00111110011010010010011011101001),
			.Kernel8(32'b00111110000001000101100100100000),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*12-1:DATA_WIDHT*11]),
			.Valid_Out(CHANNEL12_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL13 (
			.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
			.Kernel0(32'b00111110101110101011110010111011),
			.Kernel1(32'b00111111000011110100111011110011),
			.Kernel2(32'b00111110011010101100011011001100),
			.Kernel3(32'b10111111000011100001100010101110),
			.Kernel4(32'b10111110111101110001110100001111),
			.Kernel5(32'b10111110101000101101010011010111),
			.Kernel6(32'b10111110100010001010011100111000),
			.Kernel7(32'b00111110110010100111001011011101),
			.Kernel8(32'b10111110111001110101110100011010),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*13-1:DATA_WIDHT*12]),
			.Valid_Out(CHANNEL13_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL14 (
			.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
			.Kernel0(32'b00111110000110110101111100000010),
			.Kernel1(32'b10111110101010001000101000100010),
			.Kernel2(32'b00111110101110101110001011000110),
			.Kernel3(32'b00111101011101001010011001110100),
			.Kernel4(32'b00111110110001110110011010110111),
			.Kernel5(32'b10111110100000101011001110000111),
			.Kernel6(32'b00111110101011110001010110000000),
			.Kernel7(32'b00111111001000100100000101011000),
			.Kernel8(32'b00111111000001010000001111110101),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*14-1:DATA_WIDHT*13]),
			.Valid_Out(CHANNEL14_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL15 (
			.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
			.Kernel0(32'b00111110100110010110110111000001),
			.Kernel1(32'b00111100111011011100011010100101),
			.Kernel2(32'b00111110111011010110011000011011),
			.Kernel3(32'b10111110001101001101000001011110),
			.Kernel4(32'b10111111000110000000010010101010),
			.Kernel5(32'b00111101111011000010101110001100),
			.Kernel6(32'b00111111000110000111000000111011),
			.Kernel7(32'b00111110011001011010111011100110),
			.Kernel8(32'b00111110100110101111011101001100),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*15-1:DATA_WIDHT*14]),
			.Valid_Out(CHANNEL15_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL16 (
			.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
			.Kernel0(32'b10111111001001000111010011111001),
			.Kernel1(32'b10111101100101101100011111010000),
			.Kernel2(32'b10111110101111010000110100101001),
			.Kernel3(32'b00111110100000110101001011100110),
			.Kernel4(32'b00111101011011100001111110101110),
			.Kernel5(32'b10111110100011011010110001110001),
			.Kernel6(32'b00111111010001110010000100010100),
			.Kernel7(32'b00111110111010000111101000011101),
			.Kernel8(32'b00111110010010010111100101001001),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*16-1:DATA_WIDHT*15]),
			.Valid_Out(CHANNEL16_Valid_Out)
		);

endmodule