module Depthwise_Part1_Separable_64CHANNEL_Layer5  #(
    parameter DATA_WIDHT = 32, 
    parameter IMG_WIDHT = 44,
    parameter IMG_HEIGHT =44
)
(
    input [DATA_WIDHT*64-1:0] Data_In,
    input clk,
    input rst,
    input Valid_In,
    output [DATA_WIDHT*64-1:0] Data_Out,
    output Valid_Out

);
	wire CHANNEL1_Valid_Out, CHANNEL2_Valid_Out, CHANNEL3_Valid_Out, CHANNEL4_Valid_Out, CHANNEL5_Valid_Out, CHANNEL6_Valid_Out, CHANNEL7_Valid_Out, CHANNEL8_Valid_Out, CHANNEL9_Valid_Out, CHANNEL10_Valid_Out, CHANNEL11_Valid_Out, CHANNEL12_Valid_Out, CHANNEL13_Valid_Out, CHANNEL14_Valid_Out, CHANNEL15_Valid_Out, CHANNEL16_Valid_Out, CHANNEL17_Valid_Out, CHANNEL18_Valid_Out, CHANNEL19_Valid_Out, CHANNEL20_Valid_Out, CHANNEL21_Valid_Out, CHANNEL22_Valid_Out, CHANNEL23_Valid_Out, CHANNEL24_Valid_Out,CHANNEL25_Valid_Out,CHANNEL26_Valid_Out,CHANNEL27_Valid_Out,CHANNEL28_Valid_Out,CHANNEL29_Valid_Out,CHANNEL30_Valid_Out,CHANNEL31_Valid_Out,CHANNEL32_Valid_Out,CHANNEL33_Valid_Out,CHANNEL34_Valid_Out,CHANNEL35_Valid_Out,CHANNEL36_Valid_Out,CHANNEL37_Valid_Out,CHANNEL38_Valid_Out,CHANNEL39_Valid_Out,CHANNEL40_Valid_Out,CHANNEL41_Valid_Out,CHANNEL42_Valid_Out,CHANNEL43_Valid_Out,CHANNEL44_Valid_Out,CHANNEL45_Valid_Out,CHANNEL46_Valid_Out,CHANNEL47_Valid_Out,CHANNEL48_Valid_Out,CHANNEL49_Valid_Out,CHANNEL50_Valid_Out,CHANNEL51_Valid_Out,CHANNEL52_Valid_Out,CHANNEL53_Valid_Out,CHANNEL54_Valid_Out,CHANNEL55_Valid_Out,CHANNEL56_Valid_Out,CHANNEL57_Valid_Out,CHANNEL58_Valid_Out,CHANNEL59_Valid_Out,CHANNEL60_Valid_Out,CHANNEL61_Valid_Out,CHANNEL62_Valid_Out,CHANNEL63_Valid_Out,CHANNEL64_Valid_Out;

	assign Valid_Out= CHANNEL1_Valid_Out & CHANNEL2_Valid_Out & CHANNEL3_Valid_Out & CHANNEL4_Valid_Out & CHANNEL5_Valid_Out & CHANNEL6_Valid_Out & CHANNEL7_Valid_Out & CHANNEL8_Valid_Out & CHANNEL9_Valid_Out & CHANNEL10_Valid_Out & CHANNEL11_Valid_Out & CHANNEL12_Valid_Out & CHANNEL13_Valid_Out & CHANNEL14_Valid_Out & CHANNEL15_Valid_Out & CHANNEL16_Valid_Out & CHANNEL17_Valid_Out & CHANNEL18_Valid_Out & CHANNEL19_Valid_Out & CHANNEL20_Valid_Out & CHANNEL21_Valid_Out & CHANNEL22_Valid_Out& CHANNEL23_Valid_Out& CHANNEL24_Valid_Out&CHANNEL25_Valid_Out&CHANNEL26_Valid_Out&CHANNEL27_Valid_Out&CHANNEL28_Valid_Out&CHANNEL29_Valid_Out&CHANNEL30_Valid_Out&CHANNEL31_Valid_Out&CHANNEL32_Valid_Out&CHANNEL33_Valid_Out&CHANNEL34_Valid_Out&CHANNEL35_Valid_Out&CHANNEL36_Valid_Out&CHANNEL37_Valid_Out&CHANNEL38_Valid_Out&CHANNEL39_Valid_Out&CHANNEL40_Valid_Out&CHANNEL41_Valid_Out&CHANNEL42_Valid_Out&CHANNEL43_Valid_Out&CHANNEL44_Valid_Out&CHANNEL45_Valid_Out&CHANNEL46_Valid_Out&CHANNEL47_Valid_Out&CHANNEL48_Valid_Out&CHANNEL49_Valid_Out&CHANNEL50_Valid_Out&CHANNEL51_Valid_Out&CHANNEL52_Valid_Out&CHANNEL53_Valid_Out&CHANNEL54_Valid_Out&CHANNEL55_Valid_Out&CHANNEL56_Valid_Out&CHANNEL57_Valid_Out&CHANNEL58_Valid_Out&CHANNEL59_Valid_Out&CHANNEL60_Valid_Out&CHANNEL61_Valid_Out&CHANNEL62_Valid_Out&CHANNEL63_Valid_Out&CHANNEL64_Valid_Out;

	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL1 (
			.Data_In(Data_In[DATA_WIDHT-1:0]),
			.Kernel0(32'b10111110010011011000101100101101),
			.Kernel1(32'b00111110111011110001001111111100),
			.Kernel2(32'b10111110100010000110010110111000),
			.Kernel3(32'b10111100101101001111100111111001),
			.Kernel4(32'b10111111011001110000000011010010),
			.Kernel5(32'b10111110010000010111011011000001),
			.Kernel6(32'b10111100101010100111000101011100),
			.Kernel7(32'b00111111000101011110011111101010),
			.Kernel8(32'b00111111000001000100001010010000),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT-1:0]),
			.Valid_Out(CHANNEL1_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL2 (
			.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
			.Kernel0(32'b10111110001000101010110110001110),
			.Kernel1(32'b00111110100110011000110000000001),
			.Kernel2(32'b00111110110010111101011011001011),
			.Kernel3(32'b00111111000111111110001000011000),
			.Kernel4(32'b00111110000010000100010001000111),
			.Kernel5(32'b00111110110000001011000111111011),
			.Kernel6(32'b00111110011101100000111000101101),
			.Kernel7(32'b00111101010000010101000100001001),
			.Kernel8(32'b10111110100011100011111000011111),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*2-1:DATA_WIDHT]),
			.Valid_Out(CHANNEL2_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL3 (
			.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
			.Kernel0(32'b00111101000001001010100111110001),
			.Kernel1(32'b10111110111100111010100000001111),
			.Kernel2(32'b10111111001000000001001111011011),
			.Kernel3(32'b10111110100000000110100111001000),
			.Kernel4(32'b10111101101100100000110110100001),
			.Kernel5(32'b10111110101010101101001101000011),
			.Kernel6(32'b00111101111111100011010100100010),
			.Kernel7(32'b00111111000101010011011100000101),
			.Kernel8(32'b00111110100010111101011101001111),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*3-1:DATA_WIDHT*2]),
			.Valid_Out(CHANNEL3_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL4 (
			.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
			.Kernel0(32'b10111100100111100101101011101000),
			.Kernel1(32'b10111110110101010110111111100111),
			.Kernel2(32'b00111100110001011001110010111100),
			.Kernel3(32'b00111111001000000101001011001010),
			.Kernel4(32'b00111110111000000011101100101110),
			.Kernel5(32'b00111110111010111010000100001000),
			.Kernel6(32'b00111110110010101010000110110111),
			.Kernel7(32'b00111101100110100001111101011100),
			.Kernel8(32'b00111111000000101011011000011001),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*4-1:DATA_WIDHT*3]),
			.Valid_Out(CHANNEL4_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL5 (
			.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
			.Kernel0(32'b00111111000000100001101000111100),
			.Kernel1(32'b10111110100000100010100001000101),
			.Kernel2(32'b10111110010000001001001011110000),
			.Kernel3(32'b00111110101001100111010110100001),
			.Kernel4(32'b10111111000001111100010011000000),
			.Kernel5(32'b10111110110110101001111010011001),
			.Kernel6(32'b00111111001011010001111001111000),
			.Kernel7(32'b00111110000010101100111100000110),
			.Kernel8(32'b00111110110100101000000001000000),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*5-1:DATA_WIDHT*4]),
			.Valid_Out(CHANNEL5_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL6 (
			.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
			.Kernel0(32'b10111101101100001011010001011001),
			.Kernel1(32'b10111110000011110010101111001010),
			.Kernel2(32'b10111101101111101110111101010001),
			.Kernel3(32'b00111110010101011000101011101100),
			.Kernel4(32'b00111110100011000100110100100111),
			.Kernel5(32'b10111101101010110110001001100100),
			.Kernel6(32'b10111111001000110111110000101110),
			.Kernel7(32'b10111110110110001111100100110100),
			.Kernel8(32'b10111111001100101110011010011110),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*6-1:DATA_WIDHT*5]),
			.Valid_Out(CHANNEL6_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL7 (
			.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
			.Kernel0(32'b10111011101110011100001000111011),
			.Kernel1(32'b00111110111010101010111110000000),
			.Kernel2(32'b00111110111100010101010101101010),
			.Kernel3(32'b10111110101101100000110010100001),
			.Kernel4(32'b10111101000101100101000111100111),
			.Kernel5(32'b10111111001011101010001010111110),
			.Kernel6(32'b00111110110010010011101100111101),
			.Kernel7(32'b00111111001110000010001011010110),
			.Kernel8(32'b10111110010110101111001110100100),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*7-1:DATA_WIDHT*6]),
			.Valid_Out(CHANNEL7_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL8 (
			.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
			.Kernel0(32'b00111101001000011100000011000011),
			.Kernel1(32'b00111111000001110000010001110111),
			.Kernel2(32'b00111110110011101010001101010110),
			.Kernel3(32'b10111110010010000111110000001011),
			.Kernel4(32'b10111110110001111000001000100111),
			.Kernel5(32'b10111111000010110011011000110101),
			.Kernel6(32'b00111110110000110011100100000000),
			.Kernel7(32'b00111101101010100100110100111010),
			.Kernel8(32'b10111110111111000110110000010110),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*8-1:DATA_WIDHT*7]),
			.Valid_Out(CHANNEL8_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL9 (
			.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
			.Kernel0(32'b10111110010000101111101101110100),
			.Kernel1(32'b10111110101010011101100011010110),
			.Kernel2(32'b10111110111101111110001101001011),
			.Kernel3(32'b00111110111010110001010000100001),
			.Kernel4(32'b10111110110110100110101100111011),
			.Kernel5(32'b10111110000111000010111011111111),
			.Kernel6(32'b00111111001010100110011000110101),
			.Kernel7(32'b00111110100011011010001110000111),
			.Kernel8(32'b00111111001011100000110111110001),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*9-1:DATA_WIDHT*8]),
			.Valid_Out(CHANNEL9_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL10 (
			.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
			.Kernel0(32'b00111110011010000111000011100110),
			.Kernel1(32'b00111110111011101011110010001111),
			.Kernel2(32'b00111110100001011010010101111011),
			.Kernel3(32'b00111110110001001100110010101000),
			.Kernel4(32'b00111110100110100101110000101000),
			.Kernel5(32'b10111110011100100011001010101001),
			.Kernel6(32'b00111101101010110000001101011010),
			.Kernel7(32'b10111101110001010000111011011001),
			.Kernel8(32'b10111111001100111111010000111010),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*10-1:DATA_WIDHT*9]),
			.Valid_Out(CHANNEL10_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL11 (
			.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
			.Kernel0(32'b10111111000100101100001011000000),
			.Kernel1(32'b10111111010001010110011011010001),
			.Kernel2(32'b10111101111000000110011010011110),
			.Kernel3(32'b10111110001010011001101001111010),
			.Kernel4(32'b10111111000010001100100101000010),
			.Kernel5(32'b10111101101001010000010101111100),
			.Kernel6(32'b00111110011110100001101101110011),
			.Kernel7(32'b10111101000110010000100011010001),
			.Kernel8(32'b10111101010101100110010001001101),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*11-1:DATA_WIDHT*10]),
			.Valid_Out(CHANNEL11_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL12 (
			.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
			.Kernel0(32'b10111110110111100111000000100100),
			.Kernel1(32'b10111110110111010000000010100110),
			.Kernel2(32'b10111110001100000110101111010000),
			.Kernel3(32'b00111110111011001101111010011011),
			.Kernel4(32'b00111101000000011010101110101001),
			.Kernel5(32'b00111110100110011100101001010101),
			.Kernel6(32'b00111111001111101111110011001101),
			.Kernel7(32'b00111110101111101010010011101000),
			.Kernel8(32'b00111101011001010100001110101000),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*12-1:DATA_WIDHT*11]),
			.Valid_Out(CHANNEL12_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL13 (
			.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
			.Kernel0(32'b10111111000100100110000011011001),
			.Kernel1(32'b10111110101101001101100100010100),
			.Kernel2(32'b10111111001000011010000101011000),
			.Kernel3(32'b00111110000011100111001001010011),
			.Kernel4(32'b00111110010011011110000100000000),
			.Kernel5(32'b00111101110011011010101000011000),
			.Kernel6(32'b00111110111111001101001011010000),
			.Kernel7(32'b00111110000000011011001000101010),
			.Kernel8(32'b00111110100100100000001011111110),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*13-1:DATA_WIDHT*12]),
			.Valid_Out(CHANNEL13_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL14 (
			.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
			.Kernel0(32'b10111110101111111011011010111001),
			.Kernel1(32'b10111110000000001000101001011001),
			.Kernel2(32'b10111101110001001101011011000111),
			.Kernel3(32'b00111101001111111011010000100011),
			.Kernel4(32'b10111111000101001001100100111111),
			.Kernel5(32'b10111110101101110111001011011001),
			.Kernel6(32'b00111101101111000111001000011100),
			.Kernel7(32'b10111110001101001100000001110110),
			.Kernel8(32'b10111111000101001111010111100010),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*14-1:DATA_WIDHT*13]),
			.Valid_Out(CHANNEL14_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL15 (
			.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
			.Kernel0(32'b00111111001011111001101110111101),
			.Kernel1(32'b00111110011110001000110001100011),
			.Kernel2(32'b00111101111101010000100110111100),
			.Kernel3(32'b00111110111111000001101110001010),
			.Kernel4(32'b10111110111100101000000001011011),
			.Kernel5(32'b10111101100000100100100100000101),
			.Kernel6(32'b10111101100111000000101011000011),
			.Kernel7(32'b10111110000100010110110101111100),
			.Kernel8(32'b10111111001011011111111011001011),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*15-1:DATA_WIDHT*14]),
			.Valid_Out(CHANNEL15_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL16 (
			.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
			.Kernel0(32'b00111110100001011000010011010011),
			.Kernel1(32'b00111110110000011000000011111101),
			.Kernel2(32'b10111011111001100010000111010111),
			.Kernel3(32'b10111110011100110011001101101001),
			.Kernel4(32'b10111110100111110100101101001100),
			.Kernel5(32'b10111011101000001101110111110111),
			.Kernel6(32'b10111111001000111111110101110100),
			.Kernel7(32'b10111111000010110101101110010010),
			.Kernel8(32'b10111110101010111110111001100111),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*16-1:DATA_WIDHT*15]),
			.Valid_Out(CHANNEL16_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL17 (
			.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
			.Kernel0(32'b00111110101110010010011111001111),
			.Kernel1(32'b00111110111111011000100101110111),
			.Kernel2(32'b00111110001001110001000001100010),
			.Kernel3(32'b00111110100001100011000111000101),
			.Kernel4(32'b00111100011001100010010000100001),
			.Kernel5(32'b10111101001110100101100010111110),
			.Kernel6(32'b10111110111100001101010111111111),
			.Kernel7(32'b10111110110111011100101101101000),
			.Kernel8(32'b10111111010110000010100000001010),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*17-1:DATA_WIDHT*16]),
			.Valid_Out(CHANNEL17_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL18 (
			.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
			.Kernel0(32'b10111110010110010110100100101011),
			.Kernel1(32'b10111110000111001100101110001001),
			.Kernel2(32'b10111111010000011111011101011011),
			.Kernel3(32'b10111110000000010010111111110101),
			.Kernel4(32'b00111111000101111100110001111101),
			.Kernel5(32'b00111100110110101000010010000110),
			.Kernel6(32'b00111110010011110011100001110100),
			.Kernel7(32'b00111111000001111000111111001011),
			.Kernel8(32'b00111110000011100000011101100000),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*18-1:DATA_WIDHT*17]),
			.Valid_Out(CHANNEL18_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL19 (
			.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
			.Kernel0(32'b10111111010000101000101111000111),
			.Kernel1(32'b10111110010110110111010110010010),
			.Kernel2(32'b10111110010101000000111110110110),
			.Kernel3(32'b10111110111111011110001001101111),
			.Kernel4(32'b10111111000100000110110111110100),
			.Kernel5(32'b10111110010100111000101011011001),
			.Kernel6(32'b00111110100110010101010001010001),
			.Kernel7(32'b10111110000001101010001100011001),
			.Kernel8(32'b00111111000100001101110011010010),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*19-1:DATA_WIDHT*18]),
			.Valid_Out(CHANNEL19_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL20 (
			.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
			.Kernel0(32'b10111110100001110110001100111000),
			.Kernel1(32'b10111101110110001101111011011100),
			.Kernel2(32'b10111110101011000100111110000010),
			.Kernel3(32'b10111110001001110101111101110010),
			.Kernel4(32'b10111010100011010111111011001001),
			.Kernel5(32'b10111110101000001110100110101010),
			.Kernel6(32'b00111111010000111111011100111010),
			.Kernel7(32'b00111111001000111010000000001001),
			.Kernel8(32'b00111111001001011111000010010011),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*20-1:DATA_WIDHT*19]),
			.Valid_Out(CHANNEL20_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL21 (
			.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
			.Kernel0(32'b00111110111111011001110100011000),
			.Kernel1(32'b00111110000101000101100100101001),
			.Kernel2(32'b00111110100011100010000100000110),
			.Kernel3(32'b10111110110001100110101111001001),
			.Kernel4(32'b10111110101100100010000110110011),
			.Kernel5(32'b10111111010110000000110111110011),
			.Kernel6(32'b10111110110010101101101000111110),
			.Kernel7(32'b10111100001001010010111010001001),
			.Kernel8(32'b10111111001000000010010110110111),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*21-1:DATA_WIDHT*20]),
			.Valid_Out(CHANNEL21_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL22 (
			.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
			.Kernel0(32'b00111110110101001101100001101101),
			.Kernel1(32'b00111110110000001000100011000101),
			.Kernel2(32'b00111110110011100000011011000101),
			.Kernel3(32'b10111111010000110010111100000100),
			.Kernel4(32'b10111110100110111000000111100101),
			.Kernel5(32'b10111110001100010110000100111010),
			.Kernel6(32'b00111110110010011100100001010001),
			.Kernel7(32'b00111110111001110100001000011100),
			.Kernel8(32'b00111110111000100101110001011000),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*22-1:DATA_WIDHT*21]),
			.Valid_Out(CHANNEL22_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL23 (
			.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
			.Kernel0(32'b10111110111011011111100011011111),
			.Kernel1(32'b00111110011001000111001000110000),
			.Kernel2(32'b10111110100000011011000101100110),
			.Kernel3(32'b00111110101010001000001101001100),
			.Kernel4(32'b00111111001101011100011010110100),
			.Kernel5(32'b00111111001111101001111100011001),
			.Kernel6(32'b10111110010111110000111011110100),
			.Kernel7(32'b00111110000100011001111110101010),
			.Kernel8(32'b10111110100001010100011010010000),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*23-1:DATA_WIDHT*22]),
			.Valid_Out(CHANNEL23_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL24 (
			.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
			.Kernel0(32'b10111110101001010011111000111101),
			.Kernel1(32'b10111111000111111111010011100101),
			.Kernel2(32'b10111111000000010011000001100000),
			.Kernel3(32'b00111111000011110010001001001001),
			.Kernel4(32'b10111101101100110000110010110101),
			.Kernel5(32'b00111111000110010010000011000011),
			.Kernel6(32'b00111110110011011000110000111111),
			.Kernel7(32'b10111110100010100011111110010011),
			.Kernel8(32'b00111110110000110010000101001011),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*24-1:DATA_WIDHT*23]),
			.Valid_Out(CHANNEL24_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL25 (
			.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
			.Kernel0(32'b10111111001010100001000001010111),
			.Kernel1(32'b00111110011001100011100101111101),
			.Kernel2(32'b00111100110001100010100100111100),
			.Kernel3(32'b00111101110010000011110011001110),
			.Kernel4(32'b00111111001010000000001101000101),
			.Kernel5(32'b00111111000111101011100100100000),
			.Kernel6(32'b10111101000011000011100110110111),
			.Kernel7(32'b10111110001111011010101111100101),
			.Kernel8(32'b00111110000111001011110101010011),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*25-1:DATA_WIDHT*24]),
			.Valid_Out(CHANNEL25_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL26 (
			.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
			.Kernel0(32'b10111110100010111111011111110111),
			.Kernel1(32'b00111110000100101001100010011110),
			.Kernel2(32'b10111110001111111100000110001111),
			.Kernel3(32'b00111110001001011110110110010100),
			.Kernel4(32'b00111110010110110001111001110010),
			.Kernel5(32'b00111110111000010100111110010111),
			.Kernel6(32'b00111110111100100011100001100110),
			.Kernel7(32'b00111110100000111011111001100011),
			.Kernel8(32'b00111111000101100010101100110010),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*26-1:DATA_WIDHT*25]),
			.Valid_Out(CHANNEL26_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL27 (
			.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
			.Kernel0(32'b10111110010010100100111010110010),
			.Kernel1(32'b10111110111110000010111000111000),
			.Kernel2(32'b10111110000000010010010000000001),
			.Kernel3(32'b10111110100101100111111001000010),
			.Kernel4(32'b10111111000100110010001010101100),
			.Kernel5(32'b10111101111100000110010011000011),
			.Kernel6(32'b00111111001101000111110011110110),
			.Kernel7(32'b00111110111110001101001101110110),
			.Kernel8(32'b00111110110000000110001010000101),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*27-1:DATA_WIDHT*26]),
			.Valid_Out(CHANNEL27_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL28 (
			.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
			.Kernel0(32'b00111110101011110010110000010011),
			.Kernel1(32'b10111110001011000111101110011110),
			.Kernel2(32'b10111110110000101001010010001011),
			.Kernel3(32'b00111110111101110000000100101110),
			.Kernel4(32'b00111111000000011110011011011011),
			.Kernel5(32'b10111100010000101110100110101010),
			.Kernel6(32'b00111111000111100100000101001001),
			.Kernel7(32'b00111110100000100110101101110000),
			.Kernel8(32'b00111111000010111111011001110110),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*28-1:DATA_WIDHT*27]),
			.Valid_Out(CHANNEL28_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL29 (
			.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
			.Kernel0(32'b10111111000110000011111101000011),
			.Kernel1(32'b10111101010100010100011000111100),
			.Kernel2(32'b10111111001001011011100100000011),
			.Kernel3(32'b10111101110101111110001110000111),
			.Kernel4(32'b00111101111001101011110010010001),
			.Kernel5(32'b10111110001110111110011011000100),
			.Kernel6(32'b00111110000011101001000010111110),
			.Kernel7(32'b00111110010010001110001110011001),
			.Kernel8(32'b00111111010001100111001101001100),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*29-1:DATA_WIDHT*28]),
			.Valid_Out(CHANNEL29_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL30 (
			.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
			.Kernel0(32'b10111110111110001000000101010000),
			.Kernel1(32'b10111111001000101111001111101011),
			.Kernel2(32'b10111110001110111101001101100001),
			.Kernel3(32'b10111110101110000010111110010000),
			.Kernel4(32'b10111101110100101101100111111101),
			.Kernel5(32'b00111101000010011111110111010011),
			.Kernel6(32'b10111110101010000001111010100101),
			.Kernel7(32'b10111110110011011100110100101110),
			.Kernel8(32'b10111100111010101010101111000101),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*30-1:DATA_WIDHT*29]),
			.Valid_Out(CHANNEL30_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL31 (
			.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
			.Kernel0(32'b10111110111110001111010111000000),
			.Kernel1(32'b10111100111000000110111110100000),
			.Kernel2(32'b00111011000101010101000000000011),
			.Kernel3(32'b10111111001000000110001010111110),
			.Kernel4(32'b10111110001101101101100111001001),
			.Kernel5(32'b10111111001111101100110001110011),
			.Kernel6(32'b00111101101110111100000111010100),
			.Kernel7(32'b00111110101011010101010110000111),
			.Kernel8(32'b00111110000011011000110010101001),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*31-1:DATA_WIDHT*30]),
			.Valid_Out(CHANNEL31_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL32 (
			.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
			.Kernel0(32'b00111111001001111010110101010000),
			.Kernel1(32'b00111110000001111011110010010110),
			.Kernel2(32'b00111111010001011010100110110010),
			.Kernel3(32'b00111101111000110101001011110110),
			.Kernel4(32'b10111110110001000110101001100011),
			.Kernel5(32'b00111101111011100010110111100100),
			.Kernel6(32'b10111110001101000001001100001100),
			.Kernel7(32'b00111100100110111000010111111110),
			.Kernel8(32'b10111100101000001010000011001000),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*32-1:DATA_WIDHT*31]),
			.Valid_Out(CHANNEL32_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL33 (
			.Data_In(Data_In[DATA_WIDHT*33-1:DATA_WIDHT*32]),
			.Kernel0(32'b10111111000110101010101101011111),
			.Kernel1(32'b10111111000111100000010101011111),
			.Kernel2(32'b10111110111011010001001111011110),
			.Kernel3(32'b10111110111001101100111000100110),
			.Kernel4(32'b10111101100000111010011001111001),
			.Kernel5(32'b00111110100000001111000101001001),
			.Kernel6(32'b00111110101000010111001110100100),
			.Kernel7(32'b00111100011010100000100100110000),
			.Kernel8(32'b10111110101111000101011011001001),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*33-1:DATA_WIDHT*32]),
			.Valid_Out(CHANNEL33_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL34 (
			.Data_In(Data_In[DATA_WIDHT*34-1:DATA_WIDHT*33]),
			.Kernel0(32'b10111110111000110001011000110101),
			.Kernel1(32'b10111101001100101011001111001110),
			.Kernel2(32'b10111110010010110000001110010011),
			.Kernel3(32'b00111111000101010001110100010111),
			.Kernel4(32'b00111111001011110110000001010100),
			.Kernel5(32'b00111111001010100101001111100111),
			.Kernel6(32'b10111110100100111101001011010011),
			.Kernel7(32'b10111101100010011000000111111010),
			.Kernel8(32'b00111110101001100000001100111100),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*34-1:DATA_WIDHT*33]),
			.Valid_Out(CHANNEL34_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL35 (
			.Data_In(Data_In[DATA_WIDHT*35-1:DATA_WIDHT*34]),
			.Kernel0(32'b10111110101110011010001000100101),
			.Kernel1(32'b10111110111110100110101001110010),
			.Kernel2(32'b10111110111111110000001011011100),
			.Kernel3(32'b00111101110100111001000100001111),
			.Kernel4(32'b00111101111110011100111101101111),
			.Kernel5(32'b00111110101111100100111101001111),
			.Kernel6(32'b00111110111111111000100100110011),
			.Kernel7(32'b00111110100001100111010011100101),
			.Kernel8(32'b00111111000000100010101010011111),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*35-1:DATA_WIDHT*34]),
			.Valid_Out(CHANNEL35_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL36 (
			.Data_In(Data_In[DATA_WIDHT*36-1:DATA_WIDHT*35]),
			.Kernel0(32'b00111111001111010110010000011100),
			.Kernel1(32'b00111101100100101000100110010100),
			.Kernel2(32'b10111111001100111001000101011001),
			.Kernel3(32'b00111111000000010011110100110111),
			.Kernel4(32'b00111101110001111011100011101010),
			.Kernel5(32'b10111110110111001101011101000010),
			.Kernel6(32'b00111110100101110101011000110100),
			.Kernel7(32'b10111110000010000001001000010110),
			.Kernel8(32'b10111111000100100110110011100000),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*36-1:DATA_WIDHT*35]),
			.Valid_Out(CHANNEL36_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL37 (
			.Data_In(Data_In[DATA_WIDHT*37-1:DATA_WIDHT*36]),
			.Kernel0(32'b10111111000101011000001110101000),
			.Kernel1(32'b10111101111001010001011011110111),
			.Kernel2(32'b10111111001100100011111110100110),
			.Kernel3(32'b10111110111011010100110111011111),
			.Kernel4(32'b10111100110000011010010010111100),
			.Kernel5(32'b10111101011000101111000011010111),
			.Kernel6(32'b10111110101000000111100010001011),
			.Kernel7(32'b00111110100100110100111001100000),
			.Kernel8(32'b10111011110111011010110010000011),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*37-1:DATA_WIDHT*36]),
			.Valid_Out(CHANNEL37_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL38 (
			.Data_In(Data_In[DATA_WIDHT*38-1:DATA_WIDHT*37]),
			.Kernel0(32'b00111101101100011100011010111001),
			.Kernel1(32'b10111111000011011011101110101001),
			.Kernel2(32'b10111110111111000011111001010010),
			.Kernel3(32'b00111110101100110100110101001011),
			.Kernel4(32'b00111110111011100011010010110101),
			.Kernel5(32'b10111101010000110000010100011011),
			.Kernel6(32'b00111110010001011010101011000011),
			.Kernel7(32'b00111110011100100100111001010111),
			.Kernel8(32'b00111111000111100000100110100000),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*38-1:DATA_WIDHT*37]),
			.Valid_Out(CHANNEL38_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL39 (
			.Data_In(Data_In[DATA_WIDHT*39-1:DATA_WIDHT*38]),
			.Kernel0(32'b10111110000000010110111111101001),
			.Kernel1(32'b00111110001110101011011011000000),
			.Kernel2(32'b00111111000011100000100101001000),
			.Kernel3(32'b10111111001010000011001011111001),
			.Kernel4(32'b00111110000011110010011111100010),
			.Kernel5(32'b00111110011010111011011100110100),
			.Kernel6(32'b10111111001101001000110000010010),
			.Kernel7(32'b00111100010010010110100000101111),
			.Kernel8(32'b00111110101101111000110110101111),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*39-1:DATA_WIDHT*38]),
			.Valid_Out(CHANNEL39_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL40 (
			.Data_In(Data_In[DATA_WIDHT*40-1:DATA_WIDHT*39]),
			.Kernel0(32'b00111111000010001010011000100110),
			.Kernel1(32'b00111111001000001000000010111100),
			.Kernel2(32'b00111111001111011000110000111110),
			.Kernel3(32'b10111101110011010110000001110011),
			.Kernel4(32'b00111101100000001010110110010100),
			.Kernel5(32'b00111101111101001011011111000100),
			.Kernel6(32'b00111111011011000101110110010100),
			.Kernel7(32'b00111110111100100110111111100101),
			.Kernel8(32'b00111010001001001111000011011001),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*40-1:DATA_WIDHT*39]),
			.Valid_Out(CHANNEL40_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL41 (
			.Data_In(Data_In[DATA_WIDHT*41-1:DATA_WIDHT*40]),
			.Kernel0(32'b10111111001111101011011111100010),
			.Kernel1(32'b10111111010000001100010010100110),
			.Kernel2(32'b00111110110110000111101001001101),
			.Kernel3(32'b10111110111011100111111111101101),
			.Kernel4(32'b10111101100011101010010000001111),
			.Kernel5(32'b00111101011011100111111101010011),
			.Kernel6(32'b00111110001010101101101111110010),
			.Kernel7(32'b10111110001010110011110011001000),
			.Kernel8(32'b00111110101110110011011000000101),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*41-1:DATA_WIDHT*40]),
			.Valid_Out(CHANNEL41_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL42 (
			.Data_In(Data_In[DATA_WIDHT*42-1:DATA_WIDHT*41]),
			.Kernel0(32'b00111110101110110010010111001011),
			.Kernel1(32'b00111110101110011100101101000110),
			.Kernel2(32'b00111111000101110111000111011111),
			.Kernel3(32'b00111101100000000010111001101101),
			.Kernel4(32'b00111101011110010011001000100111),
			.Kernel5(32'b00111110011000001101010110100000),
			.Kernel6(32'b10111111000010010001010000110111),
			.Kernel7(32'b10111111001010010001100011010011),
			.Kernel8(32'b10111110111111001101100011101100),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*42-1:DATA_WIDHT*41]),
			.Valid_Out(CHANNEL42_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL43 (
			.Data_In(Data_In[DATA_WIDHT*43-1:DATA_WIDHT*42]),
			.Kernel0(32'b00111110101001000100010010111001),
			.Kernel1(32'b00111110101010011000000110000111),
			.Kernel2(32'b00111110111101100110110111111111),
			.Kernel3(32'b10111110001001101100001100100111),
			.Kernel4(32'b10111101001001100000100100100101),
			.Kernel5(32'b10111110001001111110001101001100),
			.Kernel6(32'b00111111000110111101011010001010),
			.Kernel7(32'b00111110101011000000111100111000),
			.Kernel8(32'b00111110101110101100101101110100),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*43-1:DATA_WIDHT*42]),
			.Valid_Out(CHANNEL43_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL44 (
			.Data_In(Data_In[DATA_WIDHT*44-1:DATA_WIDHT*43]),
			.Kernel0(32'b00111110111010011111111011101111),
			.Kernel1(32'b00111100100001111100000100000011),
			.Kernel2(32'b10111111001100110101111000101100),
			.Kernel3(32'b00111111000110101110110000001001),
			.Kernel4(32'b00111110111000011010100101110011),
			.Kernel5(32'b10111110111010110011000000101101),
			.Kernel6(32'b10111110110101001011101111101001),
			.Kernel7(32'b10111110011111111011011111010100),
			.Kernel8(32'b00111101001010110111001011110100),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*44-1:DATA_WIDHT*43]),
			.Valid_Out(CHANNEL44_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL45 (
			.Data_In(Data_In[DATA_WIDHT*45-1:DATA_WIDHT*44]),
			.Kernel0(32'b10111111010101010000010011101010),
			.Kernel1(32'b10111110101011110111101010010101),
			.Kernel2(32'b10111110011010010110001000011111),
			.Kernel3(32'b00111110111111011111101001011010),
			.Kernel4(32'b00111111000100100000011000111111),
			.Kernel5(32'b00111110101011111110000101010100),
			.Kernel6(32'b10111100110101101110110011110101),
			.Kernel7(32'b10111110011010011011110100000100),
			.Kernel8(32'b00111110101110100110111000100011),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*45-1:DATA_WIDHT*44]),
			.Valid_Out(CHANNEL45_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL46 (
			.Data_In(Data_In[DATA_WIDHT*46-1:DATA_WIDHT*45]),
			.Kernel0(32'b00111111001110101000001110001100),
			.Kernel1(32'b00111110111011001011001101111001),
			.Kernel2(32'b00111001101000001011100011100101),
			.Kernel3(32'b00111100111110011001001100011111),
			.Kernel4(32'b10111110110110110001110010001100),
			.Kernel5(32'b10111110101001101001000111010000),
			.Kernel6(32'b10111101111111000001101101100001),
			.Kernel7(32'b00111101110001011001010001011000),
			.Kernel8(32'b10111111000111001110001001111110),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*46-1:DATA_WIDHT*45]),
			.Valid_Out(CHANNEL46_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL47 (
			.Data_In(Data_In[DATA_WIDHT*47-1:DATA_WIDHT*46]),
			.Kernel0(32'b00111110111000101011001111110001),
			.Kernel1(32'b00111110110001101110110000110010),
			.Kernel2(32'b00111101110101011000001100011011),
			.Kernel3(32'b10111111001111111011111011101000),
			.Kernel4(32'b10111111000101101111100110110111),
			.Kernel5(32'b10111110111001010100111000001100),
			.Kernel6(32'b10111110011001100010100101001010),
			.Kernel7(32'b00111110011111110000111100101011),
			.Kernel8(32'b10111110010101100100101000000011),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*47-1:DATA_WIDHT*46]),
			.Valid_Out(CHANNEL47_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL48 (
			.Data_In(Data_In[DATA_WIDHT*48-1:DATA_WIDHT*47]),
			.Kernel0(32'b00111110100011011101000100011111),
			.Kernel1(32'b00111111001101001010001001011111),
			.Kernel2(32'b00111111100000110100010001011011),
			.Kernel3(32'b10111101110110111000111100001001),
			.Kernel4(32'b10111110100111110101101000000100),
			.Kernel5(32'b10111100111001001100001011101010),
			.Kernel6(32'b10111101101100011010010110100111),
			.Kernel7(32'b10111110001100100010101101110001),
			.Kernel8(32'b00111101001101010100000000001111),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*48-1:DATA_WIDHT*47]),
			.Valid_Out(CHANNEL48_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL49 (
			.Data_In(Data_In[DATA_WIDHT*49-1:DATA_WIDHT*48]),
			.Kernel0(32'b10111110100011101011100011000000),
			.Kernel1(32'b10111111001001011011100011100110),
			.Kernel2(32'b10111111010100001110111001000110),
			.Kernel3(32'b00111111000000001111100111111001),
			.Kernel4(32'b10111110011101100101000010011110),
			.Kernel5(32'b10111110110001101101001101111110),
			.Kernel6(32'b00111101100100100111111011001011),
			.Kernel7(32'b10111100011100011111100101100000),
			.Kernel8(32'b00111101101010001101101100110010),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*49-1:DATA_WIDHT*48]),
			.Valid_Out(CHANNEL49_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL50 (
			.Data_In(Data_In[DATA_WIDHT*50-1:DATA_WIDHT*49]),
			.Kernel0(32'b00111111001010110111010100111111),
			.Kernel1(32'b00111110011001110111111110010000),
			.Kernel2(32'b00111110001000011000001001000001),
			.Kernel3(32'b00111110111010111110000110001100),
			.Kernel4(32'b00111111000001110010001001110001),
			.Kernel5(32'b10111100101010101000001010010010),
			.Kernel6(32'b00111110111010010101010110111100),
			.Kernel7(32'b10111010001111101110101110001011),
			.Kernel8(32'b10111110100100000010101101111010),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*50-1:DATA_WIDHT*49]),
			.Valid_Out(CHANNEL50_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL51 (
			.Data_In(Data_In[DATA_WIDHT*51-1:DATA_WIDHT*50]),
			.Kernel0(32'b00111100110100110000001000011100),
			.Kernel1(32'b00111110111000101100011111001000),
			.Kernel2(32'b00111111001111000001111110110001),
			.Kernel3(32'b10111101010100101010011010001000),
			.Kernel4(32'b00111110100011000110001011110001),
			.Kernel5(32'b00111110001101110100111011001110),
			.Kernel6(32'b10111110110111101000001111011101),
			.Kernel7(32'b10111111000100110111101010000001),
			.Kernel8(32'b10111110100010100110110010110100),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*51-1:DATA_WIDHT*50]),
			.Valid_Out(CHANNEL51_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL52 (
			.Data_In(Data_In[DATA_WIDHT*52-1:DATA_WIDHT*51]),
			.Kernel0(32'b00111110000011111001111111111110),
			.Kernel1(32'b00111110111001100100000001000000),
			.Kernel2(32'b00111110001100111000111100100011),
			.Kernel3(32'b10111110100101001001100010001011),
			.Kernel4(32'b10111101111010000000111101001001),
			.Kernel5(32'b00111101101100111001110010010000),
			.Kernel6(32'b10111111010001001001000000000011),
			.Kernel7(32'b10111110101100110010110100001110),
			.Kernel8(32'b10111110111111011011011100111011),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*52-1:DATA_WIDHT*51]),
			.Valid_Out(CHANNEL52_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL53 (
			.Data_In(Data_In[DATA_WIDHT*53-1:DATA_WIDHT*52]),
			.Kernel0(32'b10111111010101111011010100010111),
			.Kernel1(32'b10111111000100110001101011101111),
			.Kernel2(32'b10111111001000110111101101010110),
			.Kernel3(32'b10111110000101111110110011001100),
			.Kernel4(32'b00111110101000011101111011010010),
			.Kernel5(32'b00111101001000010010010101111001),
			.Kernel6(32'b00111101101010011011100011111100),
			.Kernel7(32'b00111110001011101011011101001011),
			.Kernel8(32'b10111110000101101100101110010111),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*53-1:DATA_WIDHT*52]),
			.Valid_Out(CHANNEL53_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL54 (
			.Data_In(Data_In[DATA_WIDHT*54-1:DATA_WIDHT*53]),
			.Kernel0(32'b00111110111010000110010111100011),
			.Kernel1(32'b10111110001110001011111010111100),
			.Kernel2(32'b00111100100100000000000100110011),
			.Kernel3(32'b00111110101010011111101100110010),
			.Kernel4(32'b10111110111010001010100001111101),
			.Kernel5(32'b10111111001010011010010010110100),
			.Kernel6(32'b00111111001110101011000111000001),
			.Kernel7(32'b00111110011101111111010010111011),
			.Kernel8(32'b10111110001101110000101111000011),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*54-1:DATA_WIDHT*53]),
			.Valid_Out(CHANNEL54_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL55 (
			.Data_In(Data_In[DATA_WIDHT*55-1:DATA_WIDHT*54]),
			.Kernel0(32'b10111110001011011100110010111001),
			.Kernel1(32'b10111110100100110000101110110011),
			.Kernel2(32'b10111110010010000110111110100010),
			.Kernel3(32'b10111111000101110001100111000101),
			.Kernel4(32'b10111110101110100000111011100011),
			.Kernel5(32'b10111110110000000011010100101011),
			.Kernel6(32'b00111110111101011010100010001011),
			.Kernel7(32'b00111110101001111010111011001110),
			.Kernel8(32'b00111111000100001000000110100110),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*55-1:DATA_WIDHT*54]),
			.Valid_Out(CHANNEL55_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL56 (
			.Data_In(Data_In[DATA_WIDHT*56-1:DATA_WIDHT*55]),
			.Kernel0(32'b00111110011101001101011110001110),
			.Kernel1(32'b00111110111110101010000000100010),
			.Kernel2(32'b00111111001011011101100011100100),
			.Kernel3(32'b00111101111010001101100110100001),
			.Kernel4(32'b10111101100001000001101100000101),
			.Kernel5(32'b00111110111111101011010110111011),
			.Kernel6(32'b00111100010010010010110001001110),
			.Kernel7(32'b10111111000011011001010101000010),
			.Kernel8(32'b10111110000110011110111111101101),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*56-1:DATA_WIDHT*55]),
			.Valid_Out(CHANNEL56_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL57 (
			.Data_In(Data_In[DATA_WIDHT*57-1:DATA_WIDHT*56]),
			.Kernel0(32'b00111110111101000110010011111100),
			.Kernel1(32'b00111110001110001011010000000011),
			.Kernel2(32'b10111101110110101011001001010100),
			.Kernel3(32'b00111110111000110001000100111111),
			.Kernel4(32'b00111111000011011110001101000101),
			.Kernel5(32'b00111111001000001011110110111010),
			.Kernel6(32'b00111100111101110100001011001000),
			.Kernel7(32'b00111110001110101001010011000110),
			.Kernel8(32'b00111111001010010001010001000001),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*57-1:DATA_WIDHT*56]),
			.Valid_Out(CHANNEL57_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL58 (
			.Data_In(Data_In[DATA_WIDHT*58-1:DATA_WIDHT*57]),
			.Kernel0(32'b10111101110100011100001111000101),
			.Kernel1(32'b00111101111100111000010111101101),
			.Kernel2(32'b00111101101011110100011010011011),
			.Kernel3(32'b10111111001010011001001001000111),
			.Kernel4(32'b10111111000110011001111001100101),
			.Kernel5(32'b10111101111110101010011011100101),
			.Kernel6(32'b10111110110011111000010000110011),
			.Kernel7(32'b10111110000001100100100011101001),
			.Kernel8(32'b10111110000001101111010000110000),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*58-1:DATA_WIDHT*57]),
			.Valid_Out(CHANNEL58_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL59 (
			.Data_In(Data_In[DATA_WIDHT*59-1:DATA_WIDHT*58]),
			.Kernel0(32'b00111101111001110001001100111111),
			.Kernel1(32'b10111101110100000000101100011111),
			.Kernel2(32'b10111100101000110101011100000000),
			.Kernel3(32'b10111110011111000101010110100001),
			.Kernel4(32'b10111110011010010000001000011011),
			.Kernel5(32'b10111110111111001100010010011101),
			.Kernel6(32'b00111111001100110111111100010010),
			.Kernel7(32'b00111111000100101010100010101001),
			.Kernel8(32'b00111111000110101010000110100010),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*59-1:DATA_WIDHT*58]),
			.Valid_Out(CHANNEL59_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL60 (
			.Data_In(Data_In[DATA_WIDHT*60-1:DATA_WIDHT*59]),
			.Kernel0(32'b10111110001110010111011111000001),
			.Kernel1(32'b10111111000110101010110010111101),
			.Kernel2(32'b10111111000101010001110001111100),
			.Kernel3(32'b00111110010001110010001010011111),
			.Kernel4(32'b10111100101101011000111010110100),
			.Kernel5(32'b10111110010000001001111011111010),
			.Kernel6(32'b00111110101011110000001100000111),
			.Kernel7(32'b00111111001100110011001100100000),
			.Kernel8(32'b00111110101110011111011101010110),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*60-1:DATA_WIDHT*59]),
			.Valid_Out(CHANNEL60_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL61 (
			.Data_In(Data_In[DATA_WIDHT*61-1:DATA_WIDHT*60]),
			.Kernel0(32'b00111111000111110001001011001111),
			.Kernel1(32'b00111110101100011110010000001110),
			.Kernel2(32'b00111110101100101101111011010110),
			.Kernel3(32'b00111101100011100100001111001001),
			.Kernel4(32'b10111101010010101010010101111110),
			.Kernel5(32'b10111101001001001100010111101000),
			.Kernel6(32'b10111110110011101010101110101001),
			.Kernel7(32'b10111111001000100101100111010001),
			.Kernel8(32'b00111101101010110001001101001101),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*61-1:DATA_WIDHT*60]),
			.Valid_Out(CHANNEL61_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL62 (
			.Data_In(Data_In[DATA_WIDHT*62-1:DATA_WIDHT*61]),
			.Kernel0(32'b10111111001010000001001011011110),
			.Kernel1(32'b10111111010000101111000100000100),
			.Kernel2(32'b10111111000110100110010100110001),
			.Kernel3(32'b00111101100111111111010000110101),
			.Kernel4(32'b10111101010010111110101111011100),
			.Kernel5(32'b00111110011100111100101011110110),
			.Kernel6(32'b10111011101010110110000001101111),
			.Kernel7(32'b00111110010111011001001011100001),
			.Kernel8(32'b00111110111001001100011110110111),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*62-1:DATA_WIDHT*61]),
			.Valid_Out(CHANNEL62_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL63 (
			.Data_In(Data_In[DATA_WIDHT*63-1:DATA_WIDHT*62]),
			.Kernel0(32'b00111111001101011011010010010111),
			.Kernel1(32'b00111110100110100011000001000001),
			.Kernel2(32'b00111110001111111110111000110011),
			.Kernel3(32'b00111110101110101101100001011001),
			.Kernel4(32'b00111110010010010000111011011100),
			.Kernel5(32'b00111111000111010100101001001110),
			.Kernel6(32'b10111110101110101001000011111111),
			.Kernel7(32'b10111110010011000010001101110001),
			.Kernel8(32'b10111111001101000010100010111111),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*63-1:DATA_WIDHT*62]),
			.Valid_Out(CHANNEL63_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL64 (
			.Data_In(Data_In[DATA_WIDHT*64-1:DATA_WIDHT*63]),
			.Kernel0(32'b00111100111110011110010010100010),
			.Kernel1(32'b00111110101001110000110101001101),
			.Kernel2(32'b00111110110010010001111000010101),
			.Kernel3(32'b00111110111100011101100000000110),
			.Kernel4(32'b00111110011101001101011111011011),
			.Kernel5(32'b00111110110011111000110011011000),
			.Kernel6(32'b10111110111001100001110100111111),
			.Kernel7(32'b10111111000101100010111001100000),
			.Kernel8(32'b10111110101010110100001101000101),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*64-1:DATA_WIDHT*63]),
			.Valid_Out(CHANNEL64_Valid_Out)
		);

    
endmodule