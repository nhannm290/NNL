module Adder_64input(
    input [31:0] Data1,
    input [31:0] Data2,
    input [31:0] Data3,
    input [31:0] Data4,
    input [31:0] Data5,
    input [31:0] Data6,
    input [31:0] Data7,
    input [31:0] Data8,
    input [31:0] Data9,
    input [31:0] Data10,
    input [31:0] Data11,
    input [31:0] Data12,
    input [31:0] Data13,
    input [31:0] Data14,
    input [31:0] Data15,
    input [31:0] Data16,
    input [31:0] Data17,
    input [31:0] Data18,
    input [31:0] Data19,
    input [31:0] Data20,
    input [31:0] Data21,
    input [31:0] Data22,
    input [31:0] Data23,
    input [31:0] Data24,
    input [31:0] Data25,
    input [31:0] Data26,
    input [31:0] Data27,
    input [31:0] Data28,
    input [31:0] Data29,
    input [31:0] Data30,
    input [31:0] Data31,
    input [31:0] Data32,
    input [31:0] Data33,
    input [31:0] Data34,
    input [31:0] Data35,
    input [31:0] Data36,
    input [31:0] Data37,
    input [31:0] Data38,
    input [31:0] Data39,
    input [31:0] Data40,
    input [31:0] Data41,
    input [31:0] Data42,
    input [31:0] Data43,
    input [31:0] Data44,
    input [31:0] Data45,
    input [31:0] Data46,
    input [31:0] Data47,
    input [31:0] Data48,
    input [31:0] Data49,
    input [31:0] Data50,
    input [31:0] Data51,
    input [31:0] Data52,
    input [31:0] Data53,
    input [31:0] Data54,
    input [31:0] Data55,
    input [31:0] Data56,
    input [31:0] Data57,
    input [31:0] Data58,
    input [31:0] Data59,
    input [31:0] Data60,
    input [31:0] Data61,
    input [31:0] Data62,
    input [31:0] Data63,
    input [31:0] Data64,
    input Valid_In,
    output [31:0] Data_Out,
    output Valid_Out
);  
    wire[31:0] Data_Out1,Data_Out2;
    wire add0_Valid_Out;

    Adder_32input add0[1:0] (
        .Data1({Data1,Data17}),
        .Data2({Data2,Data18}),
        .Data3({Data3,Data19}),
        .Data4({Data4,Data20}),
        .Data5({Data5,Data21}),
        .Data6({Data6,Data22}),
        .Data7({Data7,Data23}),
        .Data8({Data8,Data24}),
        .Data9({Data9,Data25}),
        .Data10({Data10,Data26}),
        .Data11({Data11,Data27}),
        .Data12({Data12,Data28}),
        .Data13({Data13,Data29}),
        .Data14({Data14,Data30}),
        .Data15({Data15,Data31}),
        .Data16({Data16,Data32}),
        .Data17({Data33,Data49}),
        .Data18({Data34,Data50}),
        .Data19({Data35,Data51}),
        .Data20({Data36,Data52}),
        .Data21({Data37,Data53}),
        .Data22({Data38,Data54}),
        .Data23({Data39,Data55}),
        .Data24({Data40,Data56}),
        .Data25({Data41,Data57}),
        .Data26({Data42,Data58}),
        .Data27({Data43,Data59}),
        .Data28({Data44,Data60}),
        .Data29({Data45,Data61}),
        .Data30({Data46,Data62}),
        .Data31({Data47,Data63}),
        .Data32({Data48,Data64}),
        .Vadi_In(Valid_In),
        .Data_Out({Data_Out1,Data_Out2}),
        .Valid_Out(add0_Valid_Out)
    );

    FP_Adder add2 (
        .Data_A(Data_Out1), 
        .Data_B(Data_Out2),
        .Valid_In(add0_Valid_Out),
        .Mode(1'b0),
        .RMode(2'b0),
        .Data_Out(Data_Out),
        .Valid_Out(Valid_Out)
    );
    
endmodule