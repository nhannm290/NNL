module Depthwise_Part1_Separable_32CHANNEL_Layer5  #(
    parameter DATA_WIDHT = 32, 
    parameter IMG_WIDHT = 44,
    parameter IMG_HEIGHT =44
)
(
    input [DATA_WIDHT*32-1:0] Data_In,
    input clk,
    input rst,
    input Valid_In,
    output [DATA_WIDHT*32-1:0] Data_Out,
    output Valid_Out

);

	wire CHANNEL1_Valid_Out, CHANNEL2_Valid_Out, CHANNEL3_Valid_Out, CHANNEL4_Valid_Out, CHANNEL5_Valid_Out, CHANNEL6_Valid_Out, CHANNEL7_Valid_Out, CHANNEL8_Valid_Out, CHANNEL9_Valid_Out, CHANNEL10_Valid_Out, CHANNEL11_Valid_Out, CHANNEL12_Valid_Out, CHANNEL13_Valid_Out, CHANNEL14_Valid_Out, CHANNEL15_Valid_Out, CHANNEL16_Valid_Out, CHANNEL17_Valid_Out, CHANNEL18_Valid_Out, CHANNEL19_Valid_Out, CHANNEL20_Valid_Out, CHANNEL21_Valid_Out, CHANNEL22_Valid_Out, CHANNEL23_Valid_Out, CHANNEL24_Valid_Out,CHANNEL25_Valid_Out,CHANNEL26_Valid_Out,CHANNEL27_Valid_Out,CHANNEL28_Valid_Out,CHANNEL29_Valid_Out,CHANNEL30_Valid_Out,CHANNEL31_Valid_Out,CHANNEL32_Valid_Out;

	assign Valid_Out= CHANNEL1_Valid_Out & CHANNEL2_Valid_Out & CHANNEL3_Valid_Out & CHANNEL4_Valid_Out & CHANNEL5_Valid_Out & CHANNEL6_Valid_Out & CHANNEL7_Valid_Out & CHANNEL8_Valid_Out & CHANNEL9_Valid_Out & CHANNEL10_Valid_Out & CHANNEL11_Valid_Out & CHANNEL12_Valid_Out & CHANNEL13_Valid_Out & CHANNEL14_Valid_Out & CHANNEL15_Valid_Out & CHANNEL16_Valid_Out & CHANNEL17_Valid_Out & CHANNEL18_Valid_Out & CHANNEL19_Valid_Out & CHANNEL20_Valid_Out & CHANNEL21_Valid_Out & CHANNEL22_Valid_Out& CHANNEL23_Valid_Out& CHANNEL24_Valid_Out&CHANNEL25_Valid_Out&CHANNEL26_Valid_Out&CHANNEL27_Valid_Out&CHANNEL28_Valid_Out&CHANNEL29_Valid_Out&CHANNEL30_Valid_Out&CHANNEL31_Valid_Out&CHANNEL32_Valid_Out;


	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL1 (
			.Data_In(Data_In[DATA_WIDHT-1:0]),
			.Kernel0(32'b10111101010011101100101011100011),
			.Kernel1(32'b00111110011110000011100110010100),
			.Kernel2(32'b10111110101010011000010101010011),
			.Kernel3(32'b00111100001000000110110011011000),
			.Kernel4(32'b00111101111100011100110011100100),
			.Kernel5(32'b00111110000000110010001000101110),
			.Kernel6(32'b00111110110000100101010111111110),
			.Kernel7(32'b00111111000001010001010000110000),
			.Kernel8(32'b00111111000111010001011001110011),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT-1:0]),
			.Valid_Out(CHANNEL1_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL2 (
			.Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
			.Kernel0(32'b00111110111110100110110110011000),
			.Kernel1(32'b00111110000101010000000000110011),
			.Kernel2(32'b00111110100100101011110111001001),
			.Kernel3(32'b10111110100100000111010100001110),
			.Kernel4(32'b10111101100000001000010000011000),
			.Kernel5(32'b10111111000010101011010111101001),
			.Kernel6(32'b00111110001001000011011010001101),
			.Kernel7(32'b10111111001000011000010000001011),
			.Kernel8(32'b10111111000101010001010001110001),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*2-1:DATA_WIDHT]),
			.Valid_Out(CHANNEL2_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL3 (
			.Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
			.Kernel0(32'b00111110111011010110111011010110),
			.Kernel1(32'b00111101110100011111011100000100),
			.Kernel2(32'b00111111000111100011000011000010),
			.Kernel3(32'b00111111001000101101100000000011),
			.Kernel4(32'b00111101100110111101010001000000),
			.Kernel5(32'b00111110001100011111000100010100),
			.Kernel6(32'b10111110101100111101011001101010),
			.Kernel7(32'b10111110110000110111100100110000),
			.Kernel8(32'b10111110111100101110111100100110),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*3-1:DATA_WIDHT*2]),
			.Valid_Out(CHANNEL3_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL4 (
			.Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
			.Kernel0(32'b10111111001111011011101000101101),
			.Kernel1(32'b10111110100101001111100111001111),
			.Kernel2(32'b10111111000011100110101001000001),
			.Kernel3(32'b00111101111010000000001110101010),
			.Kernel4(32'b10111110100011110100000100110100),
			.Kernel5(32'b10111110010101000111100100100111),
			.Kernel6(32'b10111110101100110000110111000010),
			.Kernel7(32'b10111110001111111101011010101000),
			.Kernel8(32'b10111110100101010111011010100011),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*4-1:DATA_WIDHT*3]),
			.Valid_Out(CHANNEL4_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL5 (
			.Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
			.Kernel0(32'b10111110010011010000100011110111),
			.Kernel1(32'b00111101100100011100000010100110),
			.Kernel2(32'b10111101100010010111111000011110),
			.Kernel3(32'b10111111000000110011011010110100),
			.Kernel4(32'b10111111000101010011011001100100),
			.Kernel5(32'b10111110110110110010011101001010),
			.Kernel6(32'b00111111000000111100100101011001),
			.Kernel7(32'b00111111010101100000110011010010),
			.Kernel8(32'b00111110110100011100101000100001),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*5-1:DATA_WIDHT*4]),
			.Valid_Out(CHANNEL5_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL6 (
			.Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
			.Kernel0(32'b10111101001010110011010110001001),
			.Kernel1(32'b10111110000100010000011000010101),
			.Kernel2(32'b00111110100001010010110110011000),
			.Kernel3(32'b10111110011110100100101101111110),
			.Kernel4(32'b00111100101111101101101000010000),
			.Kernel5(32'b10111110000101010111010111111100),
			.Kernel6(32'b10111111001101110101010010101000),
			.Kernel7(32'b10111110110010111000100100100110),
			.Kernel8(32'b10111111000110000100001100110011),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*6-1:DATA_WIDHT*5]),
			.Valid_Out(CHANNEL6_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL7 (
			.Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
			.Kernel0(32'b00111111000110011011001010100110),
			.Kernel1(32'b00111110101000000100000101010010),
			.Kernel2(32'b00111111011000111000110000010000),
			.Kernel3(32'b00111110011001011010001010010110),
			.Kernel4(32'b10111100010110100110000001010010),
			.Kernel5(32'b10111110101100000001001011111110),
			.Kernel6(32'b10111111000001110011001101101100),
			.Kernel7(32'b10111111000011101000001001001100),
			.Kernel8(32'b10111101101111111100100001101111),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*7-1:DATA_WIDHT*6]),
			.Valid_Out(CHANNEL7_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL8 (
			.Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
			.Kernel0(32'b10111110100100000011111011111100),
			.Kernel1(32'b10111111000100010010110110101110),
			.Kernel2(32'b10111110100101000010000110001000),
			.Kernel3(32'b10111110011011000000110101111010),
			.Kernel4(32'b10111110111101001000011001011010),
			.Kernel5(32'b10111110011001000110111011101001),
			.Kernel6(32'b00111110001010011111101000101000),
			.Kernel7(32'b00111110010000111100001101111010),
			.Kernel8(32'b00111110101111011010000100001001),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*8-1:DATA_WIDHT*7]),
			.Valid_Out(CHANNEL8_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL9 (
			.Data_In(Data_In[DATA_WIDHT*9-1:DATA_WIDHT*8]),
			.Kernel0(32'b10111111010011010001100110100011),
			.Kernel1(32'b10111111001000001101111111010001),
			.Kernel2(32'b10111111000100011000110101110101),
			.Kernel3(32'b00111110011001111101110110000011),
			.Kernel4(32'b10111110100011110000000000100011),
			.Kernel5(32'b10111100111011001010010111001000),
			.Kernel6(32'b00111110100001000011010101100111),
			.Kernel7(32'b00111110111110000101100001000111),
			.Kernel8(32'b10111101100010100000000101100000),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*9-1:DATA_WIDHT*8]),
			.Valid_Out(CHANNEL9_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL10 (
			.Data_In(Data_In[DATA_WIDHT*10-1:DATA_WIDHT*9]),
			.Kernel0(32'b10111110011011111111101011111101),
			.Kernel1(32'b10111110110111111111011000100010),
			.Kernel2(32'b00111111010001001111001011110001),
			.Kernel3(32'b10111111000110001110011001111001),
			.Kernel4(32'b10111110110100101011001111010000),
			.Kernel5(32'b00111110011000110011000111100010),
			.Kernel6(32'b10111110111010011101011010011011),
			.Kernel7(32'b00111101011110001100011001111011),
			.Kernel8(32'b00111110010101111001101010110010),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*10-1:DATA_WIDHT*9]),
			.Valid_Out(CHANNEL10_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL11 (
			.Data_In(Data_In[DATA_WIDHT*11-1:DATA_WIDHT*10]),
			.Kernel0(32'b10111110110010000011011001001101),
			.Kernel1(32'b10111110011111110100101110000111),
			.Kernel2(32'b10111101111101011010011001001011),
			.Kernel3(32'b10111110100001010001000101100001),
			.Kernel4(32'b10111111000100111001111001001011),
			.Kernel5(32'b10111110101001000001010100100011),
			.Kernel6(32'b00111110011000100110011101110010),
			.Kernel7(32'b00111110101001110110010101010011),
			.Kernel8(32'b00111111000100100010010110000110),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*11-1:DATA_WIDHT*10]),
			.Valid_Out(CHANNEL11_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL12 (
			.Data_In(Data_In[DATA_WIDHT*12-1:DATA_WIDHT*11]),
			.Kernel0(32'b00111111001101001111101111011110),
			.Kernel1(32'b00111111001000100000101110011011),
			.Kernel2(32'b00111110000011110110000111111011),
			.Kernel3(32'b10111110000110010011011110000101),
			.Kernel4(32'b00111110000101000101110001101000),
			.Kernel5(32'b10111100001110010011111111110110),
			.Kernel6(32'b10111110110110011101101001100001),
			.Kernel7(32'b10111111000110110110100110111011),
			.Kernel8(32'b10111111001100110001001111110100),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*12-1:DATA_WIDHT*11]),
			.Valid_Out(CHANNEL12_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL13 (
			.Data_In(Data_In[DATA_WIDHT*13-1:DATA_WIDHT*12]),
			.Kernel0(32'b00111101000010111111100001011110),
			.Kernel1(32'b00111101101111100000001101100110),
			.Kernel2(32'b10111011111101000110110011000001),
			.Kernel3(32'b00111110100111110110010000100011),
			.Kernel4(32'b10111101010000000110100110111000),
			.Kernel5(32'b10111110101000001011011011100111),
			.Kernel6(32'b00111111001100001011101011100110),
			.Kernel7(32'b00111111000111101010011010100110),
			.Kernel8(32'b10111100000011001100101010111110),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*13-1:DATA_WIDHT*12]),
			.Valid_Out(CHANNEL13_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL14 (
			.Data_In(Data_In[DATA_WIDHT*14-1:DATA_WIDHT*13]),
			.Kernel0(32'b10111100101011000000000101111011),
			.Kernel1(32'b00111110010100001101100000111000),
			.Kernel2(32'b10111100001101100001110110111010),
			.Kernel3(32'b00111111000110011001011001010101),
			.Kernel4(32'b00111110111000111110010001100101),
			.Kernel5(32'b00111111000011110010111010101001),
			.Kernel6(32'b00111111000101111101011011111101),
			.Kernel7(32'b10111110001011010110001000101100),
			.Kernel8(32'b00111110100011000011001010001011),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*14-1:DATA_WIDHT*13]),
			.Valid_Out(CHANNEL14_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL15 (
			.Data_In(Data_In[DATA_WIDHT*15-1:DATA_WIDHT*14]),
			.Kernel0(32'b00111110101000000011001010011000),
			.Kernel1(32'b00111110101010111000110110000010),
			.Kernel2(32'b00111111001100110011100010110110),
			.Kernel3(32'b10111110011100101010111001011101),
			.Kernel4(32'b00111110000000000010011101110000),
			.Kernel5(32'b00111111000010101110011001011011),
			.Kernel6(32'b10111110000111101011110110111001),
			.Kernel7(32'b10111110100001100001111010111011),
			.Kernel8(32'b00111110001000111100011000101001),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*15-1:DATA_WIDHT*14]),
			.Valid_Out(CHANNEL15_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL16 (
			.Data_In(Data_In[DATA_WIDHT*16-1:DATA_WIDHT*15]),
			.Kernel0(32'b10111111000111010011011110100111),
			.Kernel1(32'b10111110110110000111101101100111),
			.Kernel2(32'b10111110000111010111110111100101),
			.Kernel3(32'b10111101100000111100000101101110),
			.Kernel4(32'b00111110000001100111011110010100),
			.Kernel5(32'b10111110000001010010101110001100),
			.Kernel6(32'b00111110110001100011011101100111),
			.Kernel7(32'b00111110100000100011110100001100),
			.Kernel8(32'b00111111001010010010000000100001),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*16-1:DATA_WIDHT*15]),
			.Valid_Out(CHANNEL16_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL17 (
			.Data_In(Data_In[DATA_WIDHT*17-1:DATA_WIDHT*16]),
			.Kernel0(32'b00111111000110100011110100000010),
			.Kernel1(32'b00111111010000101011101010101001),
			.Kernel2(32'b00111111000010011111111011110011),
			.Kernel3(32'b00111110100000101001010110101001),
			.Kernel4(32'b10111110100011111010100110000100),
			.Kernel5(32'b10111110100001110010111101000001),
			.Kernel6(32'b10111110100111001000101100010101),
			.Kernel7(32'b10111110111111101010000001001110),
			.Kernel8(32'b10111110110011010010111000100001),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*17-1:DATA_WIDHT*16]),
			.Valid_Out(CHANNEL17_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL18 (
			.Data_In(Data_In[DATA_WIDHT*18-1:DATA_WIDHT*17]),
			.Kernel0(32'b00111111010000101000101111001011),
			.Kernel1(32'b00111110101010011011110101010100),
			.Kernel2(32'b00111111001101110110010010011010),
			.Kernel3(32'b00111100110101111011110111001111),
			.Kernel4(32'b10111110001010100000011011111100),
			.Kernel5(32'b00111100001010100000010011110101),
			.Kernel6(32'b10111111000110101110001100110100),
			.Kernel7(32'b10111110101110011100011101001101),
			.Kernel8(32'b10111110011111010101101110001010),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*18-1:DATA_WIDHT*17]),
			.Valid_Out(CHANNEL18_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL19 (
			.Data_In(Data_In[DATA_WIDHT*19-1:DATA_WIDHT*18]),
			.Kernel0(32'b00111110110111110011001111001110),
			.Kernel1(32'b00111110111000111101000101000000),
			.Kernel2(32'b00111100110010000100101101110010),
			.Kernel3(32'b10111101111001010001011110010000),
			.Kernel4(32'b00111110001001111100011001000101),
			.Kernel5(32'b00111110110111010001011001100101),
			.Kernel6(32'b10111111000010011010001111100001),
			.Kernel7(32'b10111110111100110100101001011101),
			.Kernel8(32'b10111110010110100100010010010000),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*19-1:DATA_WIDHT*18]),
			.Valid_Out(CHANNEL19_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL20 (
			.Data_In(Data_In[DATA_WIDHT*20-1:DATA_WIDHT*19]),
			.Kernel0(32'b00111110101111101011000100111111),
			.Kernel1(32'b10111110001010100110011000001110),
			.Kernel2(32'b10111110100001010110011010111011),
			.Kernel3(32'b00111110110000000000101011000001),
			.Kernel4(32'b10111110001011010100101010011001),
			.Kernel5(32'b10111111011000000010010111000001),
			.Kernel6(32'b00111110111110110101010100111011),
			.Kernel7(32'b10111110100100111101011111011100),
			.Kernel8(32'b00111110001111100011111011011111),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*20-1:DATA_WIDHT*19]),
			.Valid_Out(CHANNEL20_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL21 (
			.Data_In(Data_In[DATA_WIDHT*21-1:DATA_WIDHT*20]),
			.Kernel0(32'b00111101110010101010110110000110),
			.Kernel1(32'b00111111000100110011111111010111),
			.Kernel2(32'b00111110111001001011111101100010),
			.Kernel3(32'b10111111000111001100011011111101),
			.Kernel4(32'b10111100111100010011011011010100),
			.Kernel5(32'b00111110001011001101000100100000),
			.Kernel6(32'b10111110011000010011010100101001),
			.Kernel7(32'b10111110001110001101111111000011),
			.Kernel8(32'b00111110101000110001001101100000),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*21-1:DATA_WIDHT*20]),
			.Valid_Out(CHANNEL21_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL22 (
			.Data_In(Data_In[DATA_WIDHT*22-1:DATA_WIDHT*21]),
			.Kernel0(32'b00111011111111010010011010001001),
			.Kernel1(32'b10111111000010111101000011100011),
			.Kernel2(32'b10111110001111110010100011010100),
			.Kernel3(32'b00111110011110001011000001111010),
			.Kernel4(32'b10111101100111001010000011111100),
			.Kernel5(32'b10111101111100100111101000101100),
			.Kernel6(32'b00111111001000010010000111110011),
			.Kernel7(32'b00111110111111111111101000100100),
			.Kernel8(32'b00111111000101011010000001100000),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*22-1:DATA_WIDHT*21]),
			.Valid_Out(CHANNEL22_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL23 (
			.Data_In(Data_In[DATA_WIDHT*23-1:DATA_WIDHT*22]),
			.Kernel0(32'b10111111001101011001011111101101),
			.Kernel1(32'b10111111001010110110110111001101),
			.Kernel2(32'b10111110100111111100101110110001),
			.Kernel3(32'b00111111001101110011001110011011),
			.Kernel4(32'b00111110101011100010001100111001),
			.Kernel5(32'b00111110011101100111011100010011),
			.Kernel6(32'b10111101101111000101011011000110),
			.Kernel7(32'b10111110000110011000100111010010),
			.Kernel8(32'b00111110010000101110100000111110),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*23-1:DATA_WIDHT*22]),
			.Valid_Out(CHANNEL23_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL24 (
			.Data_In(Data_In[DATA_WIDHT*24-1:DATA_WIDHT*23]),
			.Kernel0(32'b00111101101110010100110100111000),
			.Kernel1(32'b10111110010100001100101110100101),
			.Kernel2(32'b00111110011110001100000011100110),
			.Kernel3(32'b10111110001110010001111101001010),
			.Kernel4(32'b00111110110010100010010011110110),
			.Kernel5(32'b00111110100001001101101111101101),
			.Kernel6(32'b10111110101110001111111111101100),
			.Kernel7(32'b10111110110100000000110010011101),
			.Kernel8(32'b10111111011001100110100001001000),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*24-1:DATA_WIDHT*23]),
			.Valid_Out(CHANNEL24_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL25 (
			.Data_In(Data_In[DATA_WIDHT*25-1:DATA_WIDHT*24]),
			.Kernel0(32'b00111110100100111001101000001110),
			.Kernel1(32'b00111101111000101001100111011100),
			.Kernel2(32'b00111101110010011101001111111110),
			.Kernel3(32'b00111110000100101000111110111111),
			.Kernel4(32'b10111100101000011101010101001000),
			.Kernel5(32'b00111110100010000101010011101000),
			.Kernel6(32'b10111111100001101100111010111010),
			.Kernel7(32'b10111111000001001101000011000000),
			.Kernel8(32'b10111101001010000010101100110110),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*25-1:DATA_WIDHT*24]),
			.Valid_Out(CHANNEL25_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL26 (
			.Data_In(Data_In[DATA_WIDHT*26-1:DATA_WIDHT*25]),
			.Kernel0(32'b10111110101110000100111110100010),
			.Kernel1(32'b00111110001101011111000000110110),
			.Kernel2(32'b10111110101000111011000101100101),
			.Kernel3(32'b00111111000001100000110010100010),
			.Kernel4(32'b10111110010101011010101100110100),
			.Kernel5(32'b00111110011001101101100000101001),
			.Kernel6(32'b00111111000110010110111110111100),
			.Kernel7(32'b00111111000010000001100111001110),
			.Kernel8(32'b00111110100000111110100000010101),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*26-1:DATA_WIDHT*25]),
			.Valid_Out(CHANNEL26_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL27 (
			.Data_In(Data_In[DATA_WIDHT*27-1:DATA_WIDHT*26]),
			.Kernel0(32'b10111111001000100100111111011000),
			.Kernel1(32'b10111110100001010101001101101000),
			.Kernel2(32'b10111110100001100011101100000111),
			.Kernel3(32'b10111010111011011111000111111100),
			.Kernel4(32'b00111111000001111000110100110001),
			.Kernel5(32'b10111101011011110010010111000011),
			.Kernel6(32'b10111110100100101011011000000010),
			.Kernel7(32'b00111110111110010001001100001111),
			.Kernel8(32'b00111111000111101101100010001110),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*27-1:DATA_WIDHT*26]),
			.Valid_Out(CHANNEL27_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL28 (
			.Data_In(Data_In[DATA_WIDHT*28-1:DATA_WIDHT*27]),
			.Kernel0(32'b00111111000101100011100100010000),
			.Kernel1(32'b00111110111110100100000110000101),
			.Kernel2(32'b10111110110111111110000011110010),
			.Kernel3(32'b10111101111011110100011100011001),
			.Kernel4(32'b10111110110011011111110001011101),
			.Kernel5(32'b10111110100100101100110010111010),
			.Kernel6(32'b10111110010001001110111101001100),
			.Kernel7(32'b10111110000101011110011111111110),
			.Kernel8(32'b10111110101100100000101110000110),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*28-1:DATA_WIDHT*27]),
			.Valid_Out(CHANNEL28_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL29 (
			.Data_In(Data_In[DATA_WIDHT*29-1:DATA_WIDHT*28]),
			.Kernel0(32'b10111110100110100001001100010111),
			.Kernel1(32'b10111110111001011000110100110101),
			.Kernel2(32'b10111111001100100000010110001110),
			.Kernel3(32'b10111110001000101111111110110001),
			.Kernel4(32'b10111100110001111011110001001110),
			.Kernel5(32'b10111110100001001010101100001010),
			.Kernel6(32'b10111110111101110010101111011100),
			.Kernel7(32'b00111110011011101110011001001000),
			.Kernel8(32'b00111101110100010110111110011010),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*29-1:DATA_WIDHT*28]),
			.Valid_Out(CHANNEL29_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL30 (
			.Data_In(Data_In[DATA_WIDHT*30-1:DATA_WIDHT*29]),
			.Kernel0(32'b00111110001000111100111111110100),
			.Kernel1(32'b10111110000011011010000001000000),
			.Kernel2(32'b00111101111101111000000100010011),
			.Kernel3(32'b10111110011100110001000011111110),
			.Kernel4(32'b00111110110111101100101010111010),
			.Kernel5(32'b00111110011101100111110010111001),
			.Kernel6(32'b10111111001010011110000011001001),
			.Kernel7(32'b10111111010100011111100001010100),
			.Kernel8(32'b10111110100010010110000110110000),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*30-1:DATA_WIDHT*29]),
			.Valid_Out(CHANNEL30_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL31 (
			.Data_In(Data_In[DATA_WIDHT*31-1:DATA_WIDHT*30]),
			.Kernel0(32'b00111111000001101001110111001101),
			.Kernel1(32'b00111110011100000010110100101101),
			.Kernel2(32'b00111111000110001101101010110100),
			.Kernel3(32'b10111111000000011111101110010000),
			.Kernel4(32'b10111110101100001101111110110100),
			.Kernel5(32'b10111110111100110111010101111011),
			.Kernel6(32'b10111110011110010011101100010111),
			.Kernel7(32'b00111100010111001111010000001000),
			.Kernel8(32'b10111100111000111101110100100000),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*31-1:DATA_WIDHT*30]),
			.Valid_Out(CHANNEL31_Valid_Out)
		);
	Convolution2D_3x3_stride_1x1_padding_1x1 #(
		.IMG_WIDHT(IMG_WIDHT),
		.IMG_HEIGHT(IMG_HEIGHT)
	)
		CHANNEL32 (
			.Data_In(Data_In[DATA_WIDHT*32-1:DATA_WIDHT*31]),
			.Kernel0(32'b10111101110101101000100111101111),
			.Kernel1(32'b10111110011010011000100010001001),
			.Kernel2(32'b00111110011010010010111101110011),
			.Kernel3(32'b00111111000011000000010010010100),
			.Kernel4(32'b00111110111010110110110000100101),
			.Kernel5(32'b00111110101001101011110101111000),
			.Kernel6(32'b00111110010111011110100111010001),
			.Kernel7(32'b00111110100110000001101100001001),
			.Kernel8(32'b00111111000101101011011100100111),
			.Valid_In(Valid_In),
			.clk(clk),
			.rst(rst),
			.Data_Out(Data_Out[DATA_WIDHT*32-1:DATA_WIDHT*31]),
			.Valid_Out(CHANNEL32_Valid_Out)
		);

    
endmodule